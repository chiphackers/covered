module covered_top;

initial $covered_sim( "cov.cdd", top );

endmodule
