module main;

reg a = 1'b0;

endmodule
