module covered_top;

initial $covered_sim( top );

endmodule
