module main;

integer i, j;

initial begin
	i = 10 + 5 + 1 + 134;
	j = 10 + 5 + -1 + -134;
end

initial begin
        $dumpfile( "add1.vcd" );
        $dumpvars( 0, main );
        #10;
        $finish;
end

endmodule

/* HEADER
GROUPS add1 iv vcs vcd lxt
SIM    add1 iv vcd  : iverilog add1.v; ./a.out                             : add1.vcd
SIM    add1 vcs vcd : vcs add1.v;      ./simv                              : add1.vcd
SCORE  add1.vcd     : -t main -vcd add1.vcd -v add1.v -o add1.cdd          : add1.cdd
REPORT add1.cdd     : -d v -o add1.rpt add1.cdd                            : add1.rpt
*/

/* OUTPUT add1.cdd
5 1 * 6 0 0 0 0
3 0 main main add1.v 1 17
2 1 6 120014 1 0 20008 0 0 32 64 14 40 0 0 0 0 0 0
2 2 6 e000e 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 3 6 a000a 1 0 20008 0 0 32 64 11 0 0 0 0 0 0 0
2 4 6 50006 1 0 20008 0 0 32 64 44 0 0 0 0 0 0 0
2 5 6 5000a 1 6 20208 3 4 32 0 aa aa aa aa aa aa aa aa
2 6 6 5000e 1 6 20208 2 5 32 0 aa aa aa aa aa aa aa aa
2 7 6 50014 1 6 20208 1 6 32 0 aa aa aa aa aa aa aa aa
2 8 6 10001 0 1 400 0 0 i
2 9 6 10014 1 37 100a 7 8
2 10 7 140016 1 0 20008 0 0 32 64 14 40 0 0 0 0 0 0
2 11 7 130013 1 4d 20008 10 0 32 64 aa aa aa aa aa aa aa aa
2 12 7 f000f 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 13 7 e000e 1 4d 20008 12 0 32 64 aa aa aa aa aa aa aa aa
2 14 7 a000a 1 0 20008 0 0 32 64 11 0 0 0 0 0 0 0
2 15 7 50006 1 0 20008 0 0 32 64 44 0 0 0 0 0 0 0
2 16 7 5000a 1 6 20208 14 15 32 0 aa aa aa aa aa aa aa aa
2 17 7 5000f 1 6 20208 13 16 32 0 aa aa aa aa aa aa aa aa
2 18 7 50016 1 6 20208 11 17 32 0 aa aa aa aa aa aa aa aa
2 19 7 10001 0 1 400 0 0 j
2 20 7 10016 1 37 a 18 19
1 i 0 3 30008 32 112 aa aa aa aa aa aa aa aa
1 j 0 3 3000b 32 112 aa aa aa aa aa aa aa aa
4 20 0 0
4 9 20 20
*/

/* OUTPUT add1.rpt
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : add1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    add1.v                     2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    add1.v                     0/    0/    0      100%             0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              add1.v                             16/   0/  16      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    add1.v                    0/   0/   0      100%            0/   0/   0      100%


*/
