module main;

initial begin
	$dumpfile( "err2.1.vcd" );
	$dumpvars( 0, main );
end

endmodule
