module main;

parameter A = 0,
          B = 1,
          C = 2;
parameter STATE_A = (1 << A),
          STATE_B = (1 << B),
          STATE_C = (1 << C);

reg               clock;
reg [C:A]         st;
reg [C:A]         next_st;
reg [((8*8)-1):0] str;

reg  b, c, d, e, f;

always @(st or b or c or d or e or f)
  begin
   next_st = st;
   case( 1'b1 )
     st[A] :
       begin
        str = "A_STATE";
        if( b )
          next_st = STATE_B;
       end
     st[B] :
       begin
        str = "B_STATE";
        next_st = STATE_C;
       end
     st[C] :
       begin
        str = "C_STATE";
        if( c || (d && (e == f)) )
          next_st = STATE_A;
       end
   endcase
  end

always @(posedge clock) st <= next_st;
      
initial begin
	$dumpfile( "case4.vcd" );
	$dumpvars( 0, main );
	st = 3'b001;
	b  = 1'b0;
	c  = 1'b0;
	d  = 1'b0;
	e  = 1'b0;
	f  = 1'b0;
	#5;
	b  = 1'b1;
	#20;
	d  = 1'b1;
	#10;
	$finish;
end

initial begin
	clock = 1'b0;
	forever #(2) clock = ~clock;
end

endmodule

/* HEADER
GROUPS case4 all iv vcs vcd lxt
SIM    case4 all iv vcd  : iverilog case4.v; ./a.out                             : case4.vcd
SIM    case4 all iv lxt  : iverilog case4.v; ./a.out -lxt2; mv case4.vcd case4.lxt : case4.lxt
SIM    case4 all vcs vcd : vcs case4.v; ./simv                                   : case4.vcd
SCORE  case4.vcd     : -t main -vcd case4.vcd -o case4.cdd -v case4.v : case4.cdd
SCORE  case4.lxt     : -t main -lxt case4.lxt -o case4.cdd -v case4.v : case4.cdd
REPORT case4.cdd 1   : -d v -o case4.rptM case4.cdd                         : case4.rptM
REPORT case4.cdd 2   : -d v -w -o case4.rptWM case4.cdd                     : case4.rptWM
REPORT case4.cdd 3   : -d v -i -o case4.rptI case4.cdd                      : case4.rptI
REPORT case4.cdd 4   : -d v -w -i -o case4.rptWI case4.cdd                  : case4.rptWI
*/

/* OUTPUT case4.cdd
5 1 * 6 0 0 0 0
3 0 main main case4.v 1 65
2 1 19 d000e 6 1 8 0 0 st
2 2 19 30009 0 1 400 0 0 next_st
2 3 19 3000e 8 37 a 1 2
2 4 23 e0016 1 0 20008 0 0 56 4 11 10 10 11 1 10 10 11 5 11 55 11 1 10
2 5 23 8000a 0 1 400 0 0 str
2 6 23 80016 3 37 a 4 5
2 7 25 14001a 1 32 8 0 0 #STATE_B
2 8 25 a0010 0 1 400 0 0 next_st
2 9 25 a001a 2 37 600a 7 8
2 10 24 c000c 2 1 c 0 0 b
2 11 24 8000e 3 39 400e 10 0
2 12 29 e0016 1 0 20008 0 0 56 4 11 10 10 11 1 10 10 11 5 11 55 11 4 10
2 13 29 8000a 0 1 400 0 0 str
2 14 29 80016 2 37 a 12 13
2 15 30 120018 1 32 8 0 0 #STATE_C
2 16 30 8000e 0 1 400 0 0 next_st
2 17 30 80018 2 37 600a 15 16
2 18 34 e0016 1 0 20008 0 0 56 4 11 10 10 11 1 10 10 11 5 11 55 11 5 10
2 19 34 8000a 0 1 400 0 0 str
2 20 34 80016 3 37 a 18 19
2 21 36 14001a 1 32 8 0 0 #STATE_A
2 22 36 a0010 0 1 400 0 0 next_st
2 23 36 a001a 2 37 600a 21 22
2 24 35 1d001d 1 1 4 0 0 f
2 25 35 180018 1 1 4 0 0 e
2 26 35 18001d 1 11 20048 24 25 1 0 2
2 27 35 120012 2 1 c 0 0 d
2 28 35 12001e 2 18 2028c 26 27 1 0 102
2 29 35 c000c 1 1 4 0 0 c
2 30 35 c001f 2 17 200cc 28 29 1 0 102
2 31 35 80021 3 39 400e 30 0
2 32 32 80008 2 32 8 0 0 #C
2 33 32 50009 2 23 8 0 32 st
2 34 20 9000c 10 0 2000a 0 0 1 1 1
2 35 32 0 3 2d 2420a 33 34 1 0 2
2 36 27 80008 4 32 8 0 0 #B
2 37 27 50009 4 23 c 0 36 st
2 38 27 0 5 2d 2030e 37 34 1 0 1102
2 39 21 80008 6 32 4 0 0 #A
2 40 21 50009 6 23 c 0 39 st
2 41 21 0 8 2d 2030e 40 34 1 0 1102
2 42 17 230023 1 1 4 0 0 f
2 43 17 230023 0 2a 20000 0 0 2 0 a
2 44 17 230023 1 29 20008 42 43 1 0 2
2 45 17 1e001e 1 1 4 0 0 e
2 46 17 1e001e 0 2a 20000 0 0 2 0 a
2 47 17 1e001e 1 29 20008 45 46 1 0 2
2 48 17 190019 2 1 c 0 0 d
2 49 17 190019 0 2a 20000 0 0 2 0 10a
2 50 17 190019 2 29 20008 48 49 1 0 2
2 51 17 140014 1 1 4 0 0 c
2 52 17 140014 0 2a 20000 0 0 2 0 a
2 53 17 140014 1 29 20008 51 52 1 0 2
2 54 17 f000f 2 1 c 0 0 b
2 55 17 f000f 0 2a 20000 0 0 2 0 10a
2 56 17 f000f 2 29 20008 54 55 1 0 2
2 57 17 9000a 6 1 8 0 0 st
2 58 17 9000a 0 2a 20000 0 0 4 0 77aa
2 59 17 9000a 6 29 20008 57 58 1 0 2
2 60 17 9000f 7 2b 20008 56 59 1 0 2
2 61 17 90014 7 2b 20008 53 60 1 0 2
2 62 17 90019 8 2b 20008 50 61 1 0 2
2 63 17 9001e 8 2b 20008 47 62 1 0 2
2 64 17 90023 11 2b 2100a 44 63 1 0 2
2 65 41 1e0024 7 1 18 0 0 next_st
2 66 41 180019 0 1 400 0 0 st
2 67 41 180024 9 38 602a 65 66
2 68 41 110015 13 1 c 0 0 clock
2 69 41 9000f 0 2a 20000 0 0 2 0 a
2 70 41 90015 1d 27 2100a 68 69 1 0 2
2 71 61 9000c 1 0 20004 0 0 1 1 0
2 72 61 10005 0 1 400 0 0 clock
2 73 61 1000c 1 37 1006 71 72
2 74 62 17001b 12 1 1c 0 0 clock
2 75 62 160016 12 1b 2002c 74 0 1 0 1102
2 76 62 e0012 0 1 400 0 0 clock
2 77 62 e001b 12 37 602e 75 76
2 78 62 b000b 1 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 79 62 b000b 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 80 62 9000c 27 2c 2000a 78 79 32 0 aa aa aa aa aa aa aa aa
1 #A 0 0 0 32 0 0 0 0 0 0 0 0 0
1 #B 0 0 0 32 0 1 0 0 0 0 0 0 0
1 #C 0 0 0 32 0 4 0 0 0 0 0 0 0
1 #STATE_A 0 0 0 32 0 101 0 0 0 0 0 0 0
1 #STATE_B 0 0 0 32 0 204 0 0 0 0 0 0 0
1 #STATE_C 0 0 0 32 0 410 0 0 0 0 0 0 0
1 clock 0 10 30012 1 16 1102
1 st 0 11 30012 3 0 772a
1 next_st 0 12 30012 3 16 772a
1 str 0 13 30012 64 16 aa aa aa aa aa aa aa aa aa aa aa aa 33aa aa aa aa
1 b 0 15 30005 1 0 102
1 c 0 15 30008 1 0 2
1 d 0 15 3000b 1 0 102
1 e 0 15 3000e 1 0 2
1 f 0 15 30011 1 0 2
4 23 64 64
4 31 23 64
4 20 31 31
4 35 20 64
4 17 64 64
4 14 17 17
4 38 14 35
4 9 64 64
4 11 9 64
4 6 11 11
4 41 6 38
4 3 41 41
4 64 3 0
4 67 70 70
4 70 67 0
4 77 80 80
4 80 77 0
4 73 80 80
*/

/* OUTPUT case4.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : case4.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.v                   14/    0/   14      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.v                   11/   65/   76       14%             9/   67/   76       12%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      str                       0->1: 64'h0003_0000_0000_0000
      ......................... 1->0: 64'h0003_0000_0000_0000 ...
      b                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              case4.v                            18/   7/  25       72%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             19:    next_st =  st
                              |1|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             35:    if( ( c  || ( d  && ( e  ==  f ))) )
                                        |----1-----|    
                                |---------2---------|   
                        |-------------3--------------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 2   (2/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *     

        Expression 3   (2/4)
        ^^^^^^^^^^^^^ - ||
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             41:     st <= next_st
                           |--1--|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.v                   0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT case4.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : case4.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.v                   14/    0/   14      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.v                   11/   65/   76       14%             9/   67/   76       12%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      str                       0->1: 64'h0003_0000_0000_0000
      ......................... 1->0: 64'h0003_0000_0000_0000 ...
      b                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              case4.v                            18/   7/  25       72%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             19:    next_st =  st
                              |1|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             35:    if( ( c  || ( d  && ( e  ==  f ))) )
                                        |----1-----|    
                                |---------2---------|   
                        |-------------3--------------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 2   (2/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *     

        Expression 3   (2/4)
        ^^^^^^^^^^^^^ - ||
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             41:     st <= next_st
                           |--1--|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.v                   0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT case4.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : case4.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         14/    0/   14      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         11/   65/   76       14%             9/   67/   76       12%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      str                       0->1: 64'h0003_0000_0000_0000
      ......................... 1->0: 64'h0003_0000_0000_0000 ...
      b                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            18/   7/  25       72%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             19:    next_st =  st
                              |1|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             35:    if( ( c  || ( d  && ( e  ==  f ))) )
                                        |----1-----|    
                                |---------2---------|   
                        |-------------3--------------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 2   (2/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *     

        Expression 3   (2/4)
        ^^^^^^^^^^^^^ - ||
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             41:     st <= next_st
                           |--1--|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT case4.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : case4.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         14/    0/   14      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         11/   65/   76       14%             9/   67/   76       12%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      str                       0->1: 64'h0003_0000_0000_0000
      ......................... 1->0: 64'h0003_0000_0000_0000 ...
      b                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            18/   7/  25       72%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             19:    next_st =  st
                              |1|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             35:    if( ( c  || ( d  && ( e  ==  f ))) )
                                        |----1-----|    
                                |---------2---------|   
                        |-------------3--------------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 2   (2/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *     

        Expression 3   (2/4)
        ^^^^^^^^^^^^^ - ||
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             41:     st <= next_st
                           |--1--|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
