module dummy;

endmodule
