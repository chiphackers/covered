module main;

reg always_latch;

endmodule
