module main;

reg do;

endmodule
