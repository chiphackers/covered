module main;

reg priority;

endmodule
