module main;

parameter STATE_IDLE = 1'b0,
          STATE_SEND = 1'b1;

reg            clock;
reg            reset;
reg            state;
reg  [1:0]     next_state;
wire           msg_ip;
reg            head;
reg            valid;

always @(posedge clock) state <= reset ? STATE_IDLE : next_state[1];

always @(state or head or valid)
  begin
   casez( {reset, state} )
     {1'b1, 1'b?}       :  next_state = STATE_IDLE;
     {1'b0, STATE_IDLE} :  next_state = (valid & head) ? {STATE_SEND,1'b0} : {STATE_IDLE,1'b1};
     {1'b0, STATE_SEND} :  next_state =  valid         ? {STATE_SEND,1'b0} : {STATE_IDLE,1'b1};
   endcase
  end

assign msg_ip = ~next_state[0];

initial begin
	$dumpfile( "fsm5.3.vcd" );
	$dumpvars( 0, main );
	reset = 1'b1;
	valid = 1'b0;
	head  = 1'b0;
	#20;
	reset = 1'b0;
	@(posedge clock);
        head  <= 1'b1;
        valid <= 1'b1;
	@(posedge clock);
        head  <= 1'b0;
	valid <= 1'b0;
	#20;
	$finish;
end

initial begin
	clock = 1'b0;
	forever #(1) clock = ~clock;
end

endmodule

/* HEADER
GROUPS fsm5.3 all iv vcs vcd lxt
SIM    fsm5.3 all iv vcd  : iverilog fsm5.3.v; ./a.out                             : fsm5.3.vcd
SIM    fsm5.3 all iv lxt  : iverilog fsm5.3.v; ./a.out -lxt2; mv fsm5.3.vcd fsm5.3.lxt : fsm5.3.lxt
SIM    fsm5.3 all vcs vcd : vcs fsm5.3.v; ./simv                                   : fsm5.3.vcd
SCORE  fsm5.3.vcd     : -t main -vcd fsm5.3.vcd -o fsm5.3.cdd -v fsm5.3.v -F "main={reset,state},next_state[1]" : fsm5.3.cdd
SCORE  fsm5.3.lxt     : -t main -lxt fsm5.3.lxt -o fsm5.3.cdd -v fsm5.3.v -F "main={reset,state},next_state[1]" : fsm5.3.cdd
REPORT fsm5.3.cdd 1   : -d v -o fsm5.3.rptM fsm5.3.cdd                         : fsm5.3.rptM
REPORT fsm5.3.cdd 2   : -d v -w -o fsm5.3.rptWM fsm5.3.cdd                     : fsm5.3.rptWM
REPORT fsm5.3.cdd 3   : -d v -i -o fsm5.3.rptI fsm5.3.cdd                      : fsm5.3.rptI
REPORT fsm5.3.cdd 4   : -d v -w -i -o fsm5.3.rptWI fsm5.3.cdd                  : fsm5.3.rptWI
*/

/* OUTPUT fsm5.3.cdd
5 1 * 6 0 0 0 0
3 0 main main fsm5.3.v 1 50
2 1 14 410041 5 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 2 14 360042 5 23 c 0 1 next_state
2 3 14 290032 1 32 4 0 0 #STATE_IDLE
2 4 14 210032 6 1a 200cc 2 3 32 0 11aa aa aa aa aa aa aa aa
2 5 14 210025 2 1 c 0 0 reset
2 6 14 210042 6 19 201cc 4 5 1 0 1102
2 7 14 18001c 0 1 400 0 0 state
2 8 14 180042 16 38 600e 6 7
2 9 14 110015 2c 1 c 0 0 clock
2 10 14 9000f 0 2a 20000 0 0 2 0 a
2 11 14 90015 43 27 2100a 9 10 1 0 2
2 12 19 280031 1 32 4 0 0 #STATE_IDLE
2 13 19 1b0024 0 1 400 0 0 next_state
2 14 19 1b0031 2 37 6006 12 13
2 15 20 59005c 1 0 20008 0 0 1 1 1
2 16 20 4e0057 1 32 4 0 0 #STATE_IDLE
2 17 20 4e005c 1 31 20088 15 16 33 0 aa aa aa aa aa aa aa aa 2
2 18 20 4d005d 1 26 20008 17 0 33 0 aa aa aa aa aa aa aa aa 2
2 19 20 450048 1 0 20004 0 0 1 1 0
2 20 20 3a0043 1 32 8 0 0 #STATE_SEND
2 21 20 3a0048 1 31 20108 19 20 33 0 aa aa aa aa aa aa aa aa 2
2 22 20 390049 1 26 20008 21 0 33 0 aa aa aa aa aa aa aa aa 2
2 23 20 280049 2 1a 20208 18 22 33 0 21aa aa aa aa aa aa aa aa 2
2 24 20 310034 2 1 c 0 0 head
2 25 20 29002d 2 1 c 0 0 valid
2 26 20 290034 2 8 2024c 24 25 1 0 1002
2 27 20 28005d 2 19 20288 23 26 2 0 210a
2 28 20 1b0024 0 1 400 0 0 next_state
2 29 20 1b005d 2 37 600a 27 28
2 30 21 59005c 1 0 20008 0 0 1 1 1
2 31 21 4e0057 1 32 4 0 0 #STATE_IDLE
2 32 21 4e005c 1 31 20088 30 31 33 0 aa aa aa aa aa aa aa aa 2
2 33 21 4d005d 1 26 20008 32 0 33 0 aa aa aa aa aa aa aa aa 2
2 34 21 450048 1 0 20004 0 0 1 1 0
2 35 21 3a0043 1 32 8 0 0 #STATE_SEND
2 36 21 3a0048 1 31 20108 34 35 33 0 aa aa aa aa aa aa aa aa 2
2 37 21 390049 1 26 20008 36 0 33 0 aa aa aa aa aa aa aa aa 2
2 38 21 290049 1 1a 20208 33 37 33 0 aa aa aa aa aa aa aa aa 2
2 39 21 29002d 1 1 4 0 0 valid
2 40 21 29005d 1 19 20088 38 39 2 0 a
2 41 21 1b0024 0 1 400 0 0 next_state
2 42 21 1b005d 1 37 600a 40 41
2 43 21 c0015 1 32 8 0 0 #STATE_SEND
2 44 21 60009 1 0 20004 0 0 1 1 0
2 45 21 60015 1 31 20088 43 44 33 0 aa aa aa aa aa aa aa aa 2
2 46 21 50016 1 26 20008 45 0 33 0 aa aa aa aa aa aa aa aa 2
2 47 18 120016 4 1 c 0 0 state
2 48 18 b000f 2 1 c 0 0 reset
2 49 18 b0016 5 31 201cc 47 48 2 0 310a
2 50 18 a0017 9 26 2000e 49 0 2 0 310a
2 51 21 0 1 2f 2420a 46 50 1 0 2
2 52 20 c0015 1 32 4 0 0 #STATE_IDLE
2 53 20 60009 1 0 20004 0 0 1 1 0
2 54 20 60015 1 31 20044 52 53 33 0 aa aa aa aa aa aa aa aa 2
2 55 20 50016 1 26 20004 54 0 33 0 aa aa aa aa aa aa aa aa 2
2 56 20 0 3 2f 2014e 55 50 1 0 1102
2 57 19 c000f 1 0 20000 0 0 1 1 3
2 58 19 60009 1 0 20008 0 0 1 1 1
2 59 19 6000f 1 31 20008 57 58 2 0 a
2 60 19 50010 1 26 20008 59 0 2 0 a
2 61 19 0 5 2f 2028e 60 50 1 0 1002
2 62 16 1a001e 3 1 c 0 0 valid
2 63 16 1a001e 0 2a 20000 0 0 2 0 110a
2 64 16 1a001e 3 29 20008 62 63 1 0 2
2 65 16 120015 3 1 c 0 0 head
2 66 16 120015 0 2a 20000 0 0 2 0 110a
2 67 16 120015 3 29 20008 65 66 1 0 2
2 68 16 9000d 4 1 c 0 0 state
2 69 16 9000d 0 2a 20000 0 0 2 0 110a
2 70 16 9000d 4 29 20008 68 69 1 0 2
2 71 16 90015 5 2b 20008 67 70 1 0 2
2 72 16 9001e b 2b 2100a 64 71 1 0 2
2 73 25 1c001c 6 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 74 25 11001d 6 23 c 0 73 next_state
2 75 25 100010 6 1b 2000c 74 0 1 0 1002
2 76 25 7000c 0 1 400 0 0 msg_ip
2 77 25 7001d 3 35 f00e 75 76
2 78 46 9000c 1 0 20004 0 0 1 1 0
2 79 46 10005 0 1 400 0 0 clock
2 80 46 1000c 1 37 1006 78 79
2 81 47 17001b 2b 1 1c 0 0 clock
2 82 47 160016 2b 1b 2002c 81 0 1 0 1102
2 83 47 e0012 0 1 400 0 0 clock
2 84 47 e001b 2b 37 602e 82 83
2 85 47 b000b 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 86 47 b000b 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 87 47 9000c 57 2c 2000a 85 86 32 0 aa aa aa aa aa aa aa aa
2 88 0 0 6 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 89 0 0 6 23 f00e 0 88 next_state
2 90 0 0 4 1 c 0 0 state
2 91 0 0 2 1 c 0 0 reset
2 92 0 0 5 31 201cc 90 91 2 0 310a
2 93 0 0 5 26 2f00e 92 0 2 0 310a
1 #STATE_IDLE 0 0 0 32 0 0 0 0 0 0 0 0 0
1 #STATE_SEND 0 0 0 32 0 1 0 0 0 0 0 0 0
1 clock 0 6 3000f 1 16 1102
1 reset 0 7 3000f 1 0 1002
1 state 0 8 3000f 1 0 1102
1 next_state 0 9 3000f 2 16 230a
1 msg_ip 0 10 3000f 1 0 1002
1 head 0 11 3000f 1 0 1102
1 valid 0 12 3000f 1 0 1102
4 93 93 93
4 89 89 89
4 8 11 11
4 11 8 0
4 42 72 72
4 51 42 72
4 29 72 72
4 56 29 51
4 14 72 72
4 61 14 56
4 72 61 0
4 77 77 77
4 84 87 87
4 87 84 0
4 80 87 87
6 93 89 1 01,03,03,,012141
*/

/* OUTPUT fsm5.3.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm5.3.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.3.v                   9/    0/    9      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.3.v                   6/    2/    8       75%             7/    1/    8       88%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      next_state                0->1: 2'h3
      ......................... 1->0: 2'h2 ...
      msg_ip                    0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm5.3.v                           33/   5/  38       87%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             20:    next_state = (valid & head) ? {STATE_SEND, 1'b0} : {STATE_IDLE, 1'b1}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    next_state = valid ? {STATE_SEND, 1'b0} : {STATE_IDLE, 1'b1}
                                 |-1-|                                          
                                 |----------------------2----------------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
             *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.3.v                  2/  ? /  ?        ? %            3/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state ({reset, state}), output state (next_state[1])

        Hit States

          States
          ======
          1'h0
          1'h1

        Hit State Transitions

          From State    To State  
          ==========    ==========
          1'h0       -> 1'h0      
          1'h0       -> 1'h1      
          1'h1       -> 1'h0      



*/

/* OUTPUT fsm5.3.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm5.3.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.3.v                   9/    0/    9      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.3.v                   6/    2/    8       75%             7/    1/    8       88%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      next_state                0->1: 2'h3
      ......................... 1->0: 2'h2 ...
      msg_ip                    0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm5.3.v                           33/   5/  38       87%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             20:    next_state = (valid & head) ? {STATE_SEND, 1'b0} : {STATE_IDLE, 1'b1}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    next_state = valid ? {STATE_SEND, 1'b0} : {STATE_IDLE, 1'b1}
                                 |-1-|                                          
                                 |----------------------2----------------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
             *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.3.v                  2/  ? /  ?        ? %            3/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state ({reset, state}), output state (next_state[1])

        Hit States

          States
          ======
          1'h0
          1'h1

        Hit State Transitions

          From State    To State  
          ==========    ==========
          1'h0       -> 1'h0      
          1'h0       -> 1'h1      
          1'h1       -> 1'h0      



*/

/* OUTPUT fsm5.3.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm5.3.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    0/    9      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          6/    2/    8       75%             7/    1/    8       88%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      next_state                0->1: 2'h3
      ......................... 1->0: 2'h2 ...
      msg_ip                    0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            33/   5/  38       87%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             20:    next_state = (valid & head) ? {STATE_SEND, 1'b0} : {STATE_IDLE, 1'b1}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    next_state = valid ? {STATE_SEND, 1'b0} : {STATE_IDLE, 1'b1}
                                 |-1-|                                          
                                 |----------------------2----------------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
             *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         2/  ? /  ?        ? %            3/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state ({reset, state}), output state (next_state[1])

        Hit States

          States
          ======
          1'h0
          1'h1

        Hit State Transitions

          From State    To State  
          ==========    ==========
          1'h0       -> 1'h0      
          1'h0       -> 1'h1      
          1'h1       -> 1'h0      



*/

/* OUTPUT fsm5.3.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm5.3.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    0/    9      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          6/    2/    8       75%             7/    1/    8       88%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      next_state                0->1: 2'h3
      ......................... 1->0: 2'h2 ...
      msg_ip                    0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            33/   5/  38       87%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             20:    next_state = (valid & head) ? {STATE_SEND, 1'b0} : {STATE_IDLE, 1'b1}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    next_state = valid ? {STATE_SEND, 1'b0} : {STATE_IDLE, 1'b1}
                                 |-1-|                                          
                                 |----------------------2----------------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
             *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         2/  ? /  ?        ? %            3/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state ({reset, state}), output state (next_state[1])

        Hit States

          States
          ======
          1'h0
          1'h1

        Hit State Transitions

          From State    To State  
          ==========    ==========
          1'h0       -> 1'h0      
          1'h0       -> 1'h1      
          1'h1       -> 1'h0      



*/
