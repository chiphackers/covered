module main;

reg [3:0] a;
wire      b2;

foo bar[const_func(2)-1:0] (
  .a(a)
);

assign b2 = bar[3].b | bar[2].b;

initial begin
        $dumpfile( "static_func2.1.vcd" );
        $dumpvars( 0, main );
	a = 4'h4;
	#10;
	a = 4'hb;
        #10;
        $finish;
end

function [31:0] const_func;
  input [31:0] bit_to_set;
  begin
    const_func = 0;
    const_func[bit_to_set] = 1'b1;
  end
endfunction

endmodule


module foo ( input wire a );

wire b = ~a;

endmodule

/* HEADER
GROUPS static_func2.1 all vcs vcd
SIM    static_func2.1 all vcs vcd : vcs +v2k static_func2.1.v; ./simv                                     : static_func2.1.vcd
SCORE  static_func2.1.vcd     : -t main -vcd static_func2.1.vcd -o static_func2.1.cdd -v static_func2.1.v : static_func2.1.cdd
SCORE  static_func2.1.lxt     : -t main -lxt static_func2.1.lxt -o static_func2.1.cdd -v static_func2.1.v : static_func2.1.cdd
REPORT static_func2.1.cdd 1   : -d v -o static_func2.1.rptM static_func2.1.cdd                         : static_func2.1.rptM
REPORT static_func2.1.cdd 2   : -d v -w -o static_func2.1.rptWM static_func2.1.cdd                     : static_func2.1.rptWM
REPORT static_func2.1.cdd 3   : -d v -i -o static_func2.1.rptI static_func2.1.cdd                      : static_func2.1.rptI
REPORT static_func2.1.cdd 4   : -d v -w -i -o static_func2.1.rptWI static_func2.1.cdd                  : static_func2.1.rptWI
*/

/* OUTPUT static_func2.1.cdd
5 1 * 6 0 0 0 0
3 0 main main static_func2.1.v 1 30
2 1 10 17001e 2 1 c 0 0 bar[2].b
2 2 10 c0013 2 1 c 0 0 bar[3].b
2 3 10 c001e 2 9 20188 1 2 1 0 2
2 4 10 70008 0 1 400 0 0 b2
2 5 10 7001e 1 35 f00a 3 4
1 a 0 3 3000a 4 0 4baa
1 b2 0 4 3000a 1 0 2
4 5 5 5
3 0 foo main.bar[0] static_func2.1.v 33 37
2 6 35 a000a 2 1 c 0 0 a
2 7 35 90009 2 1b 2000c 6 0 1 0 1002
2 8 35 50005 0 1 400 0 0 b
2 9 35 5000a 2 36 f00e 7 8
1 a 0 33 18 1 0 102
1 b 0 35 30005 1 0 1002
4 9 9 9
3 0 foo main.bar[1] static_func2.1.v 33 37
2 30 35 a000a 2 1 c 0 0 a
2 31 35 90009 2 1b 2000c 30 0 1 0 1002
2 32 35 50005 0 1 400 0 0 b
2 33 35 5000a 2 36 f00e 31 32
1 a 0 33 18 1 0 102
1 b 0 35 30005 1 0 1002
4 33 33 33
3 0 foo main.bar[2] static_func2.1.v 33 37
2 30 35 a000a 2 1 c 0 0 a
2 31 35 90009 2 1b 2000c 30 0 1 0 102
2 32 35 50005 0 1 400 0 0 b
2 33 35 5000a 2 36 f00e 31 32
1 a 0 33 18 1 0 1002
1 b 0 35 30005 1 0 102
4 33 33 33
3 0 foo main.bar[3] static_func2.1.v 33 37
2 30 35 a000a 2 1 c 0 0 a
2 31 35 90009 2 1b 2000c 30 0 1 0 1002
2 32 35 50005 0 1 400 0 0 b
2 33 35 5000a 2 36 f00e 31 32
1 a 0 33 18 1 0 102
1 b 0 35 30005 1 0 1002
4 33 33 33
3 2 main.const_func main.const_func static_func2.1.v 22 28
2 22 25 110011 0 0 20810 0 0 32 64 0 0 0 0 0 0 0 0
2 23 25 4000d 0 1 c00 0 0 const_func
2 24 25 40011 1 37 11826 22 23
2 25 26 1d0020 0 0 20810 0 0 1 1 1
2 26 26 f0018 0 1 c00 0 0 bit_to_set
2 27 26 40019 0 23 c00 0 26 const_func
2 28 26 40020 1 37 82a 25 27
1 const_func 0 22 50010 32 16 4aa aa aa aa aa aa aa aa
1 bit_to_set 0 23 f 32 16 aa aa aa aa aa aa aa aa
4 28 0 0
4 24 28 28
*/

/* OUTPUT static_func2.1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : static_func2.1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.1.v           1/    0/    1      100%
  foo                     static_func2.1.v           1/    0/    1      100%
  main.const_func         static_func2.1.v           2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.1.v           3/    2/    5       60%             1/    4/    5       20%
  foo                     static_func2.1.v           2/    0/    2      100%             2/    0/    2      100%
  main.const_func         static_func2.1.v           1/   63/   64        2%             0/   64/   64        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'hb
      ......................... 1->0: 4'h4 ...
      b2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Function: main.const_func, File: static_func2.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      const_func                0->1: 32'h0000_0004
      ......................... 1->0: 32'h0000_0000 ...
      bit_to_set                0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              static_func2.1.v                    2/   2/   4       50%
  foo                               static_func2.1.v                    2/   0/   2      100%
  main.const_func                   static_func2.1.v                    0/   0/   0      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    assign  b2 = (bar[3].b | bar[2].b)
                                 |---------1---------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *              *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.1.v          0/   0/   0      100%            0/   0/   0      100%
  foo                     static_func2.1.v          0/   0/   0      100%            0/   0/   0      100%
  main.const_func         static_func2.1.v          0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT static_func2.1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : static_func2.1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.1.v           1/    0/    1      100%
  foo                     static_func2.1.v           1/    0/    1      100%
  main.const_func         static_func2.1.v           2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.1.v           3/    2/    5       60%             1/    4/    5       20%
  foo                     static_func2.1.v           2/    0/    2      100%             2/    0/    2      100%
  main.const_func         static_func2.1.v           1/   63/   64        2%             0/   64/   64        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'hb
      ......................... 1->0: 4'h4 ...
      b2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Function: main.const_func, File: static_func2.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      const_func                0->1: 32'h0000_0004
      ......................... 1->0: 32'h0000_0000 ...
      bit_to_set                0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              static_func2.1.v                    2/   2/   4       50%
  foo                               static_func2.1.v                    2/   0/   2      100%
  main.const_func                   static_func2.1.v                    0/   0/   0      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    assign  b2 = (bar[3].b | bar[2].b)
                                 |---------1---------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *              *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.1.v          0/   0/   0      100%            0/   0/   0      100%
  foo                     static_func2.1.v          0/   0/   0      100%            0/   0/   0      100%
  main.const_func         static_func2.1.v          0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT static_func2.1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : static_func2.1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/    0/    1      100%
  <NA>.main.bar[0]                                   1/    0/    1      100%
  <NA>.main.bar[1]                                   1/    0/    1      100%
  <NA>.main.bar[2]                                   1/    0/    1      100%
  <NA>.main.bar[3]                                   1/    0/    1      100%
  <NA>.main.const_func                               2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          3/    2/    5       60%             1/    4/    5       20%
  <NA>.main.bar[0]                                   1/    1/    2       50%             1/    1/    2       50%
  <NA>.main.bar[1]                                   1/    1/    2       50%             1/    1/    2       50%
  <NA>.main.bar[2]                                   1/    1/    2       50%             1/    1/    2       50%
  <NA>.main.bar[3]                                   1/    1/    2       50%             1/    1/    2       50%
  <NA>.main.const_func                               1/   63/   64        2%             0/   64/   64        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'hb
      ......................... 1->0: 4'h4 ...
      b2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.1.v, Instance: <NA>.main.bar[0]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: foo, File: static_func2.1.v, Instance: <NA>.main.bar[1]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: foo, File: static_func2.1.v, Instance: <NA>.main.bar[2]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      b                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.1.v, Instance: <NA>.main.bar[3]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Function: main.const_func, File: static_func2.1.v, Instance: <NA>.main.const_func
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      const_func                0->1: 32'h0000_0004
      ......................... 1->0: 32'h0000_0000 ...
      bit_to_set                0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             2/   2/   4       50%
  <NA>.main.bar[0]                                                      2/   0/   2      100%
  <NA>.main.bar[1]                                                      2/   0/   2      100%
  <NA>.main.bar[2]                                                      2/   0/   2      100%
  <NA>.main.bar[3]                                                      2/   0/   2      100%
  <NA>.main.const_func                                                  0/   0/   0      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    assign  b2 = (bar[3].b | bar[2].b)
                                 |---------1---------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *              *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[0]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[1]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[2]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[3]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.const_func                              0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT static_func2.1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : static_func2.1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/    0/    1      100%
  <NA>.main.bar[0]                                   1/    0/    1      100%
  <NA>.main.bar[1]                                   1/    0/    1      100%
  <NA>.main.bar[2]                                   1/    0/    1      100%
  <NA>.main.bar[3]                                   1/    0/    1      100%
  <NA>.main.const_func                               2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          3/    2/    5       60%             1/    4/    5       20%
  <NA>.main.bar[0]                                   1/    1/    2       50%             1/    1/    2       50%
  <NA>.main.bar[1]                                   1/    1/    2       50%             1/    1/    2       50%
  <NA>.main.bar[2]                                   1/    1/    2       50%             1/    1/    2       50%
  <NA>.main.bar[3]                                   1/    1/    2       50%             1/    1/    2       50%
  <NA>.main.const_func                               1/   63/   64        2%             0/   64/   64        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'hb
      ......................... 1->0: 4'h4 ...
      b2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.1.v, Instance: <NA>.main.bar[0]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: foo, File: static_func2.1.v, Instance: <NA>.main.bar[1]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: foo, File: static_func2.1.v, Instance: <NA>.main.bar[2]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      b                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.1.v, Instance: <NA>.main.bar[3]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Function: main.const_func, File: static_func2.1.v, Instance: <NA>.main.const_func
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      const_func                0->1: 32'h0000_0004
      ......................... 1->0: 32'h0000_0000 ...
      bit_to_set                0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             2/   2/   4       50%
  <NA>.main.bar[0]                                                      2/   0/   2      100%
  <NA>.main.bar[1]                                                      2/   0/   2      100%
  <NA>.main.bar[2]                                                      2/   0/   2      100%
  <NA>.main.bar[3]                                                      2/   0/   2      100%
  <NA>.main.const_func                                                  0/   0/   0      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    assign  b2 = (bar[3].b | bar[2].b)
                                 |---------1---------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *              *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[0]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[1]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[2]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[3]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.const_func                              0/   0/   0      100%            0/   0/   0      100%


*/
