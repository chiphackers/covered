module main;

reg         go;
reg         a;
reg         b, c;
reg  [27:3] d;
reg         e;

always @(posedge go)
  begin
   a = (b | c) &
         ((d[27:16]==12'h0) &&
         (d[12:3] != 10'h000) &&
         (d[12:3] != 10'h001) &&
         (d[12:3] != 10'h002) &&
         (d[12:3] != 10'h003) &&
         (d[12:3] != 10'h004) &&
         (d[12:3] != 10'h005) &&
         (d[12:3] != 10'h006) &&
         (d[12:3] != 10'h007) &&
         (d[12:3] != 10'h008) &&
         (d[12:3] != 10'h009) &&
         (d[12:3] != 10'h00A) &&
         (d[12:3] != 10'h00B) &&
         (d[12:3] != 10'h00C) &&
         (d[12:3] != 10'h00D) &&
         (d[12:3] != 10'h00E) &&
         (d[12:3] != 10'h00F) &&
         (d[12:3] != 10'h010) &&
         (d[12:3] != 10'h011) &&
         (d[12:3] != 10'h012) &&
         (d[12:3] != 10'h013) &&
         (d[12:3] != 10'h014) &&
         (d[12:3] != 10'h015) &&
         (d[12:3] != 10'h016) &&
         (d[12:3] != 10'h017) &&
         (d[12:3] != 10'h018) &&
         (d[12:3] != 10'h019) &&
         (d[12:3] != 10'h01A) &&
         (d[12:3] != 10'h01B) &&
         (d[12:3] != 10'h01C) &&
         (d[12:3] != 10'h01D) &&
         (d[12:3] != 10'h01E) &&
         (d[12:3] != 10'h01F) &&
         (d[12:3] != 10'h020) &&
         (d[12:3] != 10'h021) &&
         (d[12:3] != 10'h022) &&
         (d[12:3] != 10'h023) &&
         (d[12:3] != 10'h024) &&
         (d[12:3] != 10'h025) &&
         (d[12:3] != 10'h026) &&
         (d[12:3] != 10'h027) &&
         (d[12:3] != 10'h028) &&
         (d[12:3] != 10'h029) &&
         (d[12:3] != 10'h02A) &&
         (d[12:3] != 10'h02B) &&
         (d[12:3] != 10'h02C) &&
         (d[12:3] != 10'h02D) &&
         (d[12:3] != 10'h02E) &&
         (d[12:3] != 10'h02F) &&
         (d[12:3] != 10'h030) &&
         (d[12:3] != 10'h031) &&
         (d[12:3] != 10'h032) &&
         (d[12:3] != 10'h033) &&
         (d[12:3] != 10'h034) &&
         (d[12:3] != 10'h035) &&
         (d[12:3] != 10'h036) &&
         (d[12:3] != 10'h037) &&
         (d[12:3] != 10'h038) &&
         (d[12:3] != 10'h039) &&
         (d[12:3] != 10'h03A) &&
         (d[12:3] != 10'h03B) &&
         (d[12:3] != 10'h03C) &&
         (d[12:3] != 10'h03D) &&
         (d[12:3] != 10'h03E) &&
         (d[12:3] != 10'h03F) &&
         (d[12:3] != 10'h040) &&
         (d[12:3] != 10'h041) &&
         (d[12:3] != 10'h042) &&
         (d[12:3] != 10'h043) &&
         (d[12:3] != 10'h044) &&
         (d[12:3] != 10'h045) &&
         (d[12:3] != 10'h046) &&
         (d[12:3] != 10'h047) &&
         (d[12:3] != 10'h048) &&
         (d[12:3] != 10'h049) &&
         (d[12:3] != 10'h04A) &&
         (d[12:3] != 10'h04B) &&
         (d[12:3] != 10'h04C) &&
         (d[12:3] != 10'h04D) &&
         (d[12:3] != 10'h04E) &&
         (d[12:3] != 10'h04F) &&
         (d[12:3] != 10'h050) &&
         (d[12:3] != 10'h051) &&
         (d[12:3] != 10'h052) &&
         (d[12:3] != 10'h053) &&
         (d[12:3] != 10'h054)) |
        e &
        ((d[27:16]==12'h0) &&
         (d[12:3] != 10'h000) &&
         (d[12:3] != 10'h001) &&
         (d[12:3] != 10'h002) &&
         (d[12:3] != 10'h003) &&
         (d[12:3] != 10'h004) &&
         (d[12:3] != 10'h005) &&
         (d[12:3] != 10'h006) &&
         (d[12:3] != 10'h007) &&
         (d[12:3] != 10'h008) &&
         (d[12:3] != 10'h009) &&
         (d[12:3] != 10'h00A) &&
         (d[12:3] != 10'h00B) &&
         (d[12:3] != 10'h00C) &&
         (d[12:3] != 10'h00D) &&
         (d[12:3] != 10'h00E) &&
         (d[12:3] != 10'h00F) &&
         (d[12:3] != 10'h010) &&
         (d[12:3] != 10'h011) &&
         (d[12:3] != 10'h012) &&
         (d[12:3] != 10'h013) &&
         (d[12:3] != 10'h014) &&
         (d[12:3] != 10'h015) &&
         (d[12:3] != 10'h016) &&
         (d[12:3] != 10'h017) &&
         (d[12:3] != 10'h018) &&
         (d[12:3] != 10'h019) &&
         (d[12:3] != 10'h01A) &&
         (d[12:3] != 10'h01B) &&
         (d[12:3] != 10'h01C) &&
         (d[12:3] != 10'h01D) &&
         (d[12:3] != 10'h01E) &&
         (d[12:3] != 10'h01F) &&
         (d[12:3] != 10'h020) &&
         (d[12:3] != 10'h021) &&
         (d[12:3] != 10'h022) &&
         (d[12:3] != 10'h023) &&
         (d[12:3] != 10'h024) &&
         (d[12:3] != 10'h025) &&
         (d[12:3] != 10'h026) &&
         (d[12:3] != 10'h027) &&
         (d[12:3] != 10'h028) &&
         (d[12:3] != 10'h029) &&
         (d[12:3] != 10'h02A) &&
         (d[12:3] != 10'h02B) &&
         (d[12:3] != 10'h02C) &&
         (d[12:3] != 10'h02D) &&
         (d[12:3] != 10'h02E) &&
         (d[12:3] != 10'h02F) &&
         (d[12:3] != 10'h030) &&
         (d[12:3] != 10'h031) &&
         (d[12:3] != 10'h032) &&
         (d[12:3] != 10'h033) &&
         (d[12:3] != 10'h034) &&
         (d[12:3] != 10'h035) &&
         (d[12:3] != 10'h036) &&
         (d[12:3] != 10'h037) &&
         (d[12:3] != 10'h038) &&
         (d[12:3] != 10'h039) &&
         (d[12:3] != 10'h03A) &&
         (d[12:3] != 10'h03B) &&
         (d[12:3] != 10'h03C) &&
         (d[12:3] != 10'h03D) &&
         (d[12:3] != 10'h03E) &&
         (d[12:3] != 10'h03F) &&
         (d[12:3] != 10'h040) &&
         (d[12:3] != 10'h041) &&
         (d[12:3] != 10'h042) &&
         (d[12:3] != 10'h043) &&
         (d[12:3] != 10'h044) &&
         (d[12:3] != 10'h045) &&
         (d[12:3] != 10'h046) &&
         (d[12:3] != 10'h047) &&
         (d[12:3] != 10'h048) &&
         (d[12:3] != 10'h049) &&
         (d[12:3] != 10'h04A) &&
         (d[12:3] != 10'h04B)) ;
  end

initial begin
	$dumpfile( "long_exp2.vcd" );
	$dumpvars( 0, main );
	b = 1'b0;
	c = 1'b0;
	d = 25'h0000000;
	e = 1'b0;
	#5;
	$finish;
end

endmodule
