module main (
  input wire a
);

endmodule
