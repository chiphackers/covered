/*
 Name:     comment1.v
 Author:   Trevor Williams  (phase1geo@gmail.com)
 Date:     11/02/2006
 Purpose:  Verifies that the parser properly parses a comment with a comment.
*/

/* This is a /* comment */ in a comment */

module main;

endmodule
