module main;

reg unique;

endmodule
