module main (
  output wire [1:0] foo
);

endmodule
