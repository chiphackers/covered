`define ST_STOP     3'b001
`define ST_GO       3'b010
`define ST_SLOW     3'b100

module main;

reg        clk;
reg        go;
wire [2:0] state;

fsma fsm1( clk, go, state );
fsmb fsm2( clk, go );

wire error = (state[0] & state[1]) || (state[0] & state[2]) || (state[1] & state[2]) || (state == 3'b000);

initial begin
	$dumpfile( "example.vcd" );
	$dumpvars( 0, main );
	go = 1'b0;
	repeat( 10 ) @(posedge clk);
	go = 1'b1;
	#10;
	$finish;
end

initial begin
	clk = 1'b0;
	forever #(1) clk = ~clk;
end

endmodule

module fsma( clk, go, state );

input        clk;
input        go;
output [2:0] state;

reg [2:0] next_state;
reg [2:0] state;

initial begin
	state = `ST_SLOW;
end

always @(posedge clk) state <= next_state;

(* covered_fsm, lights, is="state", os="next_state" *)
always @(state or go)
  case( state )
    `ST_STOP :  next_state = go ? `ST_GO : `ST_STOP;
    `ST_GO   :  next_state = go ? `ST_GO : `ST_SLOW;
    `ST_SLOW :  next_state = `ST_STOP;
  endcase

endmodule

module fsmb( clk, go );

input     clk;
input     go;
     
reg [2:0] next_state;
reg [2:0] state;  
     
initial begin
        state = `ST_STOP;
end     
        
always @(posedge clk) state <= next_state;
        
(* covered_fsm, lights, is="state", os="next_state",
                        trans="3'b001->3'b010",
                        trans="3'b010->3'b100",
                        trans="3'b100->3'b001" *)
always @(state or go)
  case( state )
    `ST_STOP :  next_state = go ? `ST_GO : `ST_STOP;
    `ST_GO   :  next_state = go ? `ST_GO : `ST_SLOW;
    `ST_SLOW :  next_state = `ST_STOP;
  endcase
        
endmodule

/* HEADER
GROUPS example all iv vcd lxt
SIM    example all iv vcd  : iverilog example.v; ./a.out                             : example.vcd
SIM    example all iv lxt  : iverilog example.v; ./a.out -lxt2; mv example.vcd example.lxt : example.lxt
SCORE  example.vcd     : -t main -vcd example.vcd -o example.cdd -v example.v : example.cdd
SCORE  example.lxt     : -t main -lxt example.lxt -o example.cdd -v example.v : example.cdd
REPORT example.cdd 1   : -d v -o example.rptM example.cdd                         : example.rptM
REPORT example.cdd 2   : -d v -w -o example.rptWM example.cdd                     : example.rptWM
REPORT example.cdd 3   : -d v -i -o example.rptI example.cdd                      : example.rptI
REPORT example.cdd 4   : -d v -w -i -o example.rptWI example.cdd                  : example.rptWI
*/

/* OUTPUT example.cdd
5 1 * 6 0 0 0 0
3 0 main main example.v 5 31
2 1 14 620067 1 0 20004 0 0 3 1 0
2 2 14 59005d 3 1 8 0 0 state
2 3 14 590067 4 11 20104 1 2 1 0 2
2 4 14 510051 4 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 5 14 4b0052 4 23 c 0 4 state
2 6 14 460046 4 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 7 14 400047 4 23 c 0 6 state
2 8 14 400052 4 8 201c4 5 7 1 0 2
2 9 14 380038 4 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 10 14 320039 4 23 c 0 9 state
2 11 14 2d002d 4 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 12 14 27002e 4 23 c 0 11 state
2 13 14 270039 4 8 201c4 10 12 1 0 2
2 14 14 1f001f 4 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 15 14 190020 4 23 c 0 14 state
2 16 14 140014 4 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 17 14 e0015 4 23 c 0 16 state
2 18 14 e0020 4 8 201c4 15 17 1 0 2
2 19 14 d003a 4 17 20044 13 18 1 0 2
2 20 14 d0053 4 17 20044 8 19 1 0 2
2 21 14 d0068 4 17 20044 3 20 1 0 2
2 22 14 50009 0 1 400 0 0 error
2 23 14 50068 2 36 f006 21 22
2 24 27 7000a 1 0 20004 0 0 1 1 0
2 25 27 10003 0 1 400 0 0 clk
2 26 27 1000a 1 37 1006 24 25
2 27 28 150017 1d 1 1c 0 0 clk
2 28 28 140014 1d 1b 2002c 27 0 1 0 1102
2 29 28 e0010 0 1 400 0 0 clk
2 30 28 e0017 1d 37 602e 28 29
2 31 28 b000b 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 32 28 b000b 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 33 28 9000c 3b 2c 2000a 31 32 32 0 aa aa aa aa aa aa aa aa
1 clk 0 7 3000b 1 16 1102
1 go 0 8 3000b 1 0 102
1 state 0 9 3000b 3 0 532a
1 error 0 14 30005 1 0 2
4 23 23 23
4 30 33 33
4 33 30 0
4 26 33 33
3 0 fsma main.fsm1 example.v 33 56
2 34 51 29002e 1 0 20008 0 0 3 1 1
2 35 51 200025 1 0 20008 0 0 3 1 4
2 36 51 1b0025 2 1a 20208 34 35 3 0 122a
2 37 51 1b001c 2 1 c 0 0 go
2 38 51 1b002e 2 19 20288 36 37 3 0 122a
2 39 51 e0017 0 1 400 0 0 next_state
2 40 51 e002e 2 37 600a 38 39
2 41 52 2b0030 1 0 20008 0 0 3 1 10
2 42 52 220027 1 0 20008 0 0 3 1 4
2 43 52 1d0027 1 1a 20208 41 42 3 0 2a
2 44 52 1d001e 1 1 8 0 0 go
2 45 52 1d0030 1 19 20208 43 44 3 0 2a
2 46 52 100019 0 1 400 0 0 next_state
2 47 52 100030 1 37 600a 45 46
2 48 53 1b0020 1 0 20008 0 0 3 1 1
2 49 53 e0017 0 1 400 0 0 next_state
2 50 53 e0020 1 37 600a 48 49
2 51 53 40009 1 0 20008 0 0 3 1 10
2 52 50 8000c 7 1 a 0 0 state
2 53 53 0 1 2d 2420a 51 52 1 0 2
2 54 52 40009 1 0 20008 0 0 3 1 4
2 55 52 0 2 2d 2020e 54 52 1 0 102
2 56 51 40009 1 0 20008 0 0 3 1 1
2 57 51 0 4 2d 2020e 56 52 1 0 1102
2 58 49 120013 2 1 c 0 0 go
2 59 49 120013 0 2a 20000 0 0 2 0 10a
2 60 49 120013 2 29 20008 58 59 1 0 2
2 61 49 9000d 3 1 8 0 0 state
2 62 49 9000d 0 2a 20000 0 0 4 0 53aa
2 63 49 9000d 3 29 20008 61 62 1 0 2
2 64 49 90013 9 2b 2100a 60 63 1 0 2
2 65 0 0 4 1 f00a 0 0 next_state
2 66 0 0 3 1 f00a 0 0 state
1 clk 0 35 d 1 0 1102
1 go 0 36 d 1 0 102
1 state 0 37 1000d 3 0 532a
1 next_state 0 39 3000a 3 16 122a
4 66 66 66
4 65 65 65
4 50 64 64
4 53 50 64
4 47 64 64
4 55 47 53
4 40 64 64
4 57 40 55
4 64 57 0
6 66 65 1 03,06,04,,2104210141014102
7 4 46 46
3 0 fsmb main.fsm2 example.v 58 83
2 67 78 29002e 1 0 20008 0 0 3 1 1
2 68 78 200025 1 0 20008 0 0 3 1 4
2 69 78 1b0025 2 1a 20208 67 68 3 0 122a
2 70 78 1b001c 2 1 c 0 0 go
2 71 78 1b002e 2 19 20288 69 70 3 0 122a
2 72 78 e0017 0 1 400 0 0 next_state
2 73 78 e002e 2 37 600a 71 72
2 74 79 2b0030 1 0 20008 0 0 3 1 10
2 75 79 220027 1 0 20008 0 0 3 1 4
2 76 79 1d0027 1 1a 20208 74 75 3 0 2a
2 77 79 1d001e 1 1 8 0 0 go
2 78 79 1d0030 1 19 20208 76 77 3 0 2a
2 79 79 100019 0 1 400 0 0 next_state
2 80 79 100030 1 37 600a 78 79
2 81 80 1b0020 0 0 20010 0 0 3 1 1
2 82 80 e0017 0 1 400 0 0 next_state
2 83 80 e0020 0 37 6022 81 82
2 84 80 40009 0 0 20010 0 0 3 1 10
2 85 77 8000c 4 1 a 0 0 state
2 86 80 0 0 2d 24022 84 85 1 0 2
2 87 79 40009 1 0 20008 0 0 3 1 4
2 88 79 0 1 2d 2020a 87 85 1 0 2
2 89 78 40009 1 0 20008 0 0 3 1 1
2 90 78 0 3 2d 2020e 89 85 1 0 1002
2 91 76 120013 2 1 c 0 0 go
2 92 76 120013 0 2a 20000 0 0 2 0 10a
2 93 76 120013 2 29 20008 91 92 1 0 2
2 94 76 9000d 2 1 8 0 0 state
2 95 76 9000d 0 2a 20000 0 0 4 0 12aa
2 96 76 9000d 2 29 20008 94 95 1 0 2
2 97 76 90013 7 2b 2100a 93 96 1 0 2
2 98 0 0 3 1 f00a 0 0 next_state
2 99 0 0 2 1 f00a 0 0 state
1 clk 0 60 a 1 0 1102
1 go 0 61 a 1 0 102
1 next_state 0 63 3000a 3 16 122a
1 state 0 64 3000a 3 0 122a
4 99 99 99
4 98 98 98
4 83 97 97
4 86 83 97
4 80 97 97
4 88 80 86
4 73 97 97
4 90 73 88
4 97 90 0
6 99 98 1 03,06,05,0141018002200421014102
7 4 70 70
*/

/* OUTPUT example.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : example.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    example.v                  3/    0/    3      100%
  fsma                    example.v                  4/    0/    4      100%
  fsmb                    example.v                  3/    1/    4       75%
---------------------------------------------------------------------------------------------------------------------

    Module: fsmb, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           80:    next_state = 3'b1



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    example.v                  4/    2/    6       67%             3/    3/    6       50%
  fsma                    example.v                  5/    3/    8       62%             4/    4/    8       50%
  fsmb                    example.v                  4/    4/    8       50%             3/    5/    8       38%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      state                     0->1: 3'h3
      ......................... 1->0: 3'h5 ...
      error                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: fsma, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      state                     0->1: 3'h3
      ......................... 1->0: 3'h5 ...
      next_state                0->1: 3'h2
      ......................... 1->0: 3'h1 ...

    Module: fsmb, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      next_state                0->1: 3'h2
      ......................... 1->0: 3'h1 ...
      state                     0->1: 3'h2
      ......................... 1->0: 3'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              example.v                          13/   8/  21       62%
  fsma                              example.v                           8/   4/  12       67%
  fsmb                              example.v                           8/   4/  12       67%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             14:    error = ((state[0] & state[1]) || (state[0] & state[2]) || (state[1] & state[2]) || (state == 3'b0))
                             |---------1---------|    |---------2---------|    |---------3---------|    |------4------| 
                            |--------------------------------------------5---------------------------------------------|

        Expression 1   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 2   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 3   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 4   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
             *

        Expression 5   (1/5)
        ^^^^^^^^^^^^^ - ||
         1 | 2 | 3 | 4 | All
        =1=|=1=|=1=|=1=|==0==
         *   *   *   *       


    Module: fsma, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             51:    case( state ) 
                          |-1-|   
                    3'b1 :

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             51:    next_state =  go ? 3'b10 : 3'b1
                                 |-------1--------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             52:    next_state =  go ? 3'b10 : 3'b100
                                 |1|                 
                                 |--------2---------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    


    Module: fsmb, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    case( state ) 
                          |-1-|   
                    3'b1 :

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    next_state =  go ? 3'b10 : 3'b1
                                 |-------1--------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             79:    next_state =  go ? 3'b10 : 3'b100
                                 |1|                 
                                 |--------2---------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    example.v                 0/   0/   0      100%            0/   0/   0      100%
  fsma                    example.v                 3/  ? /  ?        ? %            4/  ? /  ?        ? %
  fsmb                    example.v                 2/   1/   3       67%            3/   2/   5       60%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: example.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          3'h4
          3'h1
          3'h2

        Hit State Transitions

          From State    To State  
          ==========    ==========
          3'h4       -> 3'h1      
          3'h1       -> 3'h1      
          3'h1       -> 3'h2      
          3'h2       -> 3'h2      


    Module: fsmb, File: example.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          3'h4

        Missed State Transitions

          From State    To State  
          ==========    ==========
          3'h2       -> 3'h4      
          3'h4       -> 3'h1      



*/

/* OUTPUT example.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : example.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    example.v                  3/    0/    3      100%
  fsma                    example.v                  4/    0/    4      100%
  fsmb                    example.v                  3/    1/    4       75%
---------------------------------------------------------------------------------------------------------------------

    Module: fsmb, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           80:    next_state = 3'b1



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    example.v                  4/    2/    6       67%             3/    3/    6       50%
  fsma                    example.v                  5/    3/    8       62%             4/    4/    8       50%
  fsmb                    example.v                  4/    4/    8       50%             3/    5/    8       38%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      state                     0->1: 3'h3
      ......................... 1->0: 3'h5 ...
      error                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: fsma, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      state                     0->1: 3'h3
      ......................... 1->0: 3'h5 ...
      next_state                0->1: 3'h2
      ......................... 1->0: 3'h1 ...

    Module: fsmb, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      next_state                0->1: 3'h2
      ......................... 1->0: 3'h1 ...
      state                     0->1: 3'h2
      ......................... 1->0: 3'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              example.v                          13/   8/  21       62%
  fsma                              example.v                           8/   4/  12       67%
  fsmb                              example.v                           8/   4/  12       67%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             14:    error = ((state[0] & state[1]) || (state[0] & state[2]) || (state[1] & state[2]) || (state == 3'b0))
                             |---------1---------|    |---------2---------|    |---------3---------|    |------4------| 
                            |--------------------------------------------5---------------------------------------------|

        Expression 1   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 2   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 3   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 4   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
             *

        Expression 5   (1/5)
        ^^^^^^^^^^^^^ - ||
         1 | 2 | 3 | 4 | All
        =1=|=1=|=1=|=1=|==0==
         *   *   *   *       


    Module: fsma, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             51:    case( state ) 3'b1 :
                          |-1-|         

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             51:    next_state =  go ? 3'b10 : 3'b1
                                 |-------1--------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             52:    next_state =  go ? 3'b10 : 3'b100
                                 |1|                 
                                 |--------2---------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    


    Module: fsmb, File: example.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    case( state ) 3'b1 :
                          |-1-|         

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    next_state =  go ? 3'b10 : 3'b1
                                 |-------1--------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             79:    next_state =  go ? 3'b10 : 3'b100
                                 |1|                 
                                 |--------2---------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    example.v                 0/   0/   0      100%            0/   0/   0      100%
  fsma                    example.v                 3/  ? /  ?        ? %            4/  ? /  ?        ? %
  fsmb                    example.v                 2/   1/   3       67%            3/   2/   5       60%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: example.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          3'h4
          3'h1
          3'h2

        Hit State Transitions

          From State    To State  
          ==========    ==========
          3'h4       -> 3'h1      
          3'h1       -> 3'h1      
          3'h1       -> 3'h2      
          3'h2       -> 3'h2      


    Module: fsmb, File: example.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          3'h4

        Missed State Transitions

          From State    To State  
          ==========    ==========
          3'h2       -> 3'h4      
          3'h4       -> 3'h1      



*/

/* OUTPUT example.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : example.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          3/    0/    3      100%
  <NA>.main.fsm1                                     4/    0/    4      100%
  <NA>.main.fsm2                                     3/    1/    4       75%
---------------------------------------------------------------------------------------------------------------------

    Module: fsmb, File: example.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           80:    next_state = 3'b1



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          4/    2/    6       67%             3/    3/    6       50%
  <NA>.main.fsm1                                     5/    3/    8       62%             4/    4/    8       50%
  <NA>.main.fsm2                                     4/    4/    8       50%             3/    5/    8       38%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: example.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      state                     0->1: 3'h3
      ......................... 1->0: 3'h5 ...
      error                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: fsma, File: example.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      state                     0->1: 3'h3
      ......................... 1->0: 3'h5 ...
      next_state                0->1: 3'h2
      ......................... 1->0: 3'h1 ...

    Module: fsmb, File: example.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      next_state                0->1: 3'h2
      ......................... 1->0: 3'h1 ...
      state                     0->1: 3'h2
      ......................... 1->0: 3'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            13/   8/  21       62%
  <NA>.main.fsm1                                                        8/   4/  12       67%
  <NA>.main.fsm2                                                        8/   4/  12       67%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: example.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             14:    error = ((state[0] & state[1]) || (state[0] & state[2]) || (state[1] & state[2]) || (state == 3'b0))
                             |---------1---------|    |---------2---------|    |---------3---------|    |------4------| 
                            |--------------------------------------------5---------------------------------------------|

        Expression 1   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 2   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 3   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 4   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
             *

        Expression 5   (1/5)
        ^^^^^^^^^^^^^ - ||
         1 | 2 | 3 | 4 | All
        =1=|=1=|=1=|=1=|==0==
         *   *   *   *       


    Module: fsma, File: example.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             51:    case( state ) 
                          |-1-|   
                    3'b1 :

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             51:    next_state =  go ? 3'b10 : 3'b1
                                 |-------1--------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             52:    next_state =  go ? 3'b10 : 3'b100
                                 |1|                 
                                 |--------2---------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    


    Module: fsmb, File: example.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    case( state ) 
                          |-1-|   
                    3'b1 :

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    next_state =  go ? 3'b10 : 3'b1
                                 |-------1--------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             79:    next_state =  go ? 3'b10 : 3'b100
                                 |1|                 
                                 |--------2---------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.fsm1                                    3/  ? /  ?        ? %            4/  ? /  ?        ? %
  <NA>.main.fsm2                                    2/   1/   3       67%            3/   2/   5       60%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: example.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          3'h4
          3'h1
          3'h2

        Hit State Transitions

          From State    To State  
          ==========    ==========
          3'h4       -> 3'h1      
          3'h1       -> 3'h1      
          3'h1       -> 3'h2      
          3'h2       -> 3'h2      


    Module: fsmb, File: example.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          3'h4

        Missed State Transitions

          From State    To State  
          ==========    ==========
          3'h2       -> 3'h4      
          3'h4       -> 3'h1      



*/

/* OUTPUT example.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : example.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          3/    0/    3      100%
  <NA>.main.fsm1                                     4/    0/    4      100%
  <NA>.main.fsm2                                     3/    1/    4       75%
---------------------------------------------------------------------------------------------------------------------

    Module: fsmb, File: example.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           80:    next_state = 3'b1



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          4/    2/    6       67%             3/    3/    6       50%
  <NA>.main.fsm1                                     5/    3/    8       62%             4/    4/    8       50%
  <NA>.main.fsm2                                     4/    4/    8       50%             3/    5/    8       38%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: example.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      state                     0->1: 3'h3
      ......................... 1->0: 3'h5 ...
      error                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: fsma, File: example.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      state                     0->1: 3'h3
      ......................... 1->0: 3'h5 ...
      next_state                0->1: 3'h2
      ......................... 1->0: 3'h1 ...

    Module: fsmb, File: example.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      next_state                0->1: 3'h2
      ......................... 1->0: 3'h1 ...
      state                     0->1: 3'h2
      ......................... 1->0: 3'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            13/   8/  21       62%
  <NA>.main.fsm1                                                        8/   4/  12       67%
  <NA>.main.fsm2                                                        8/   4/  12       67%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: example.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             14:    error = ((state[0] & state[1]) || (state[0] & state[2]) || (state[1] & state[2]) || (state == 3'b0))
                             |---------1---------|    |---------2---------|    |---------3---------|    |------4------| 
                            |--------------------------------------------5---------------------------------------------|

        Expression 1   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 2   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 3   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                        *

        Expression 4   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
             *

        Expression 5   (1/5)
        ^^^^^^^^^^^^^ - ||
         1 | 2 | 3 | 4 | All
        =1=|=1=|=1=|=1=|==0==
         *   *   *   *       


    Module: fsma, File: example.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             51:    case( state ) 3'b1 :
                          |-1-|         

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             51:    next_state =  go ? 3'b10 : 3'b1
                                 |-------1--------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             52:    next_state =  go ? 3'b10 : 3'b100
                                 |1|                 
                                 |--------2---------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    


    Module: fsmb, File: example.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    case( state ) 3'b1 :
                          |-1-|         

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    next_state =  go ? 3'b10 : 3'b1
                                 |-------1--------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             79:    next_state =  go ? 3'b10 : 3'b100
                                 |1|                 
                                 |--------2---------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.fsm1                                    3/  ? /  ?        ? %            4/  ? /  ?        ? %
  <NA>.main.fsm2                                    2/   1/   3       67%            3/   2/   5       60%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: example.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          3'h4
          3'h1
          3'h2

        Hit State Transitions

          From State    To State  
          ==========    ==========
          3'h4       -> 3'h1      
          3'h1       -> 3'h1      
          3'h1       -> 3'h2      
          3'h2       -> 3'h2      


    Module: fsmb, File: example.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          3'h4

        Missed State Transitions

          From State    To State  
          ==========    ==========
          3'h2       -> 3'h4      
          3'h4       -> 3'h1      



*/
