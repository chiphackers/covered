module main;

reg	    a, b, c;
reg [2:0]   d;

wire        w0;
wire        w1, w2, w3, w4;
wire        w5;
wire        w6; 
wire        w7, w8, w9;
wire        w10, w11, w12, w13, w14, w15, w16, w17, w18, w19; 
wire        w20, w21, w22, w23, w24, w25, w26, w27;
wire [31:0] x0;
wire [31:0] x1; 
wire [31:0] x2; 
wire [31:0] x3, x4, x5, x6;
wire [1:0]  y0;
wire [1:0]  y1;
wire [1:0]  y2;

integer     i; 
integer     j, k, l;

assign w0 = 0;             // EXP_OP_NONE
assign w1 = a;             // EXP_OP_SIG  -- wrong
assign w2 = a ^ b;         // EXP_OP_XOR
assign x0 = a * b;         // EXP_OP_MULTIPLY
assign x1 = a / 1;         // EXP_OP_DIVIDE
assign x2 = a % 2;         // EXP_OP_MOD
assign x3 = a + b;         // EXP_OP_ADD
assign x4 = a - b;         // EXP_OP_SUBTRACT
assign w3 = a & b;	   // EXP_OP_AND
assign w4 = a | b;         // EXP_OP_OR
assign w5 = a ~& b;        // EXP_OP_NAND
assign w6 = a ~| b;        // EXP_OP_NOR
assign w7 = a ~^ b;        // EXP_OP_NXOR
assign w8 = a < b;         // EXP_OP_LT
assign w9 = a > b;         // EXP_OP_GT
assign x5 = a << b;        // EXP_OP_LSHIFT
assign x6 = a >> b;        // EXP_OP_RSHIFT
assign w10 = a == b;       // EXP_OP_EQ
assign w11 = a === b;      // EXP_OP_CEQ
assign w12 = a <= b;       // EXP_OP_LE
assign w13 = a >= b;       // EXP_OP_GE
assign w14 = a != b;       // EXP_OP_NE
assign w15 = a !== b;      // EXP_OP_CNE
assign w16 = a || b;       // EXP_OP_LOR
assign w17 = a && b;       // EXP_OP_LAND
assign w18 = a ? b : c;    // EXP_OP_COND/EXP_OP_COND_SEL
assign w19 = ~a;           // EXP_OP_UINV
assign w20 = &d;           // EXP_OP_UAND
assign w21 = !a;           // EXP_OP_UNOT
assign w22 = |d;           // EXP_OP_UOR
assign w23 = ^d;           // EXP_OP_UXOR
assign w24 = ~&d;          // EXP_OP_UNAND
assign w25 = ~|d;          // EXP_OP_UNOR
assign w26 = ~^d;          // EXP_OP_UNXOR
assign w27 = d[1];         // EXP_OP_SBIT_SEL
assign y0  = d[2:1];       // EXP_OP_MBIT_SEL
assign y1  = {2{a}};       // EXP_OP_EXPAND
assign y2  = {a, b};       // EXP_OP_CONCAT -- wrong

initial begin
	$dumpfile( "assign1.vcd" );
        $dumpvars( 0, main );
	for( i=0; i<2; i=i+1 )
          begin
           a = i;
           for( j=0; j<2; j=j+1 )
             begin
              b = j;
              for( k=0; k<2; k=k+1 )
                begin
                 c = k;
                 for( l=0; l<8; l=l+1 )
                   begin
                    d = l;
                    #5;
                   end
                end
             end
          end 
        a = 0;
        b = 0;
        #5;
end

endmodule

/* HEADER
GROUPS assign1 all iv vcd lxt
SIM    assign1 all iv vcd  : iverilog assign1.v; ./a.out                             : assign1.vcd
SIM    assign1 all iv lxt  : iverilog assign1.v; ./a.out -lxt2; mv assign1.vcd assign1.lxt : assign1.lxt
SCORE  assign1.vcd     : -t main -vcd assign1.vcd -o assign1.cdd -v assign1.v : assign1.cdd
SCORE  assign1.lxt     : -t main -lxt assign1.lxt -o assign1.cdd -v assign1.v : assign1.cdd
REPORT assign1.cdd 1   : -d v -o assign1.rptM assign1.cdd                         : assign1.rptM
REPORT assign1.cdd 2   : -d v -w -o assign1.rptWM assign1.cdd                     : assign1.rptWM
REPORT assign1.cdd 3   : -d v -i -o assign1.rptI assign1.cdd                      : assign1.rptI
REPORT assign1.cdd 4   : -d v -w -i -o assign1.rptWI assign1.cdd                  : assign1.rptWI
*/

/* OUTPUT assign1.cdd
5 1 * 6 0 0 0 0
3 0 main main assign1.v 1 88
2 1 24 c000c 1 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 2 24 70008 0 1 400 0 0 w0
2 3 24 7000c 1 35 f006 1 2
2 4 25 c000c 3 1 c 0 0 a
2 5 25 70008 0 1 400 0 0 w1
2 6 25 7000c 3 35 f00e 4 5
2 7 26 100010 5 1 c 0 0 b
2 8 26 c000c 3 1 c 0 0 a
2 9 26 c0010 5 2 203cc 7 8 1 0 1102
2 10 26 70008 0 1 400 0 0 w2
2 11 26 70010 3 35 f00e 9 10
2 12 27 100010 5 1 c 0 0 b
2 13 27 c000c 3 1 c 0 0 a
2 14 27 c0010 5 3 203cc 12 13 2 0 110a
2 15 27 70008 0 1 400 0 0 x0
2 16 27 70010 3 35 f00e 14 15
2 17 28 100010 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 18 28 c000c 3 1 c 0 0 a
2 19 28 c0010 4 4 2028c 17 18 32 0 11aa aa aa aa aa aa aa aa
2 20 28 70008 0 1 400 0 0 x1
2 21 28 70010 4 35 f00e 19 20
2 22 29 100010 1 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 23 29 c000c 3 1 c 0 0 a
2 24 29 c0010 4 5 2028c 22 23 32 0 11aa aa aa aa aa aa aa aa
2 25 29 70008 0 1 400 0 0 x2
2 26 29 70010 4 35 f00e 24 25
2 27 30 100010 5 1 c 0 0 b
2 28 30 c000c 3 1 c 0 0 a
2 29 30 c0010 5 6 203cc 27 28 32 0 33aa aa aa aa aa aa aa aa
2 30 30 70008 0 1 400 0 0 x3
2 31 30 70010 4 35 f00e 29 30
2 32 31 100010 5 1 c 0 0 b
2 33 31 c000c 3 1 c 0 0 a
2 34 31 c0010 5 7 203c8 32 33 32 0 33aa aa aa aa aa aa aa aa
2 35 31 70008 0 1 400 0 0 x4
2 36 31 70010 4 35 f00a 34 35
2 37 32 100010 5 1 c 0 0 b
2 38 32 c000c 3 1 c 0 0 a
2 39 32 c0010 5 8 203cc 37 38 1 0 1102
2 40 32 70008 0 1 400 0 0 w3
2 41 32 70010 3 35 f00e 39 40
2 42 33 100010 5 1 c 0 0 b
2 43 33 c000c 3 1 c 0 0 a
2 44 33 c0010 5 9 203cc 42 43 1 0 1102
2 45 33 70008 0 1 400 0 0 w4
2 46 33 70010 3 35 f00e 44 45
2 47 34 110011 5 1 c 0 0 b
2 48 34 c000c 3 1 c 0 0 a
2 49 34 c0011 5 a 203cc 47 48 1 0 1102
2 50 34 70008 0 1 400 0 0 w5
2 51 34 70011 3 35 f00e 49 50
2 52 35 110011 5 1 c 0 0 b
2 53 35 c000c 3 1 c 0 0 a
2 54 35 c0011 5 b 203cc 52 53 1 0 1102
2 55 35 70008 0 1 400 0 0 w6
2 56 35 70011 3 35 f00e 54 55
2 57 36 110011 5 1 c 0 0 b
2 58 36 c000c 3 1 c 0 0 a
2 59 36 c0011 5 c 203cc 57 58 1 0 1102
2 60 36 70008 0 1 400 0 0 w7
2 61 36 70011 3 35 f00e 59 60
2 62 37 100010 5 1 c 0 0 b
2 63 37 c000c 3 1 c 0 0 a
2 64 37 c0010 5 d 203cc 62 63 1 0 1102
2 65 37 70008 0 1 400 0 0 w8
2 66 37 70010 3 35 f00e 64 65
2 67 38 100010 5 1 c 0 0 b
2 68 38 c000c 3 1 c 0 0 a
2 69 38 c0010 5 e 203cc 67 68 1 0 1102
2 70 38 70008 0 1 400 0 0 w9
2 71 38 70010 3 35 f00e 69 70
2 72 39 110011 5 1 c 0 0 b
2 73 39 c000c 3 1 c 0 0 a
2 74 39 c0011 5 f 203cc 72 73 32 0 11aa aa aa aa aa aa aa aa
2 75 39 70008 0 1 400 0 0 x5
2 76 39 70011 3 35 f00e 74 75
2 77 40 110011 5 1 c 0 0 b
2 78 40 c000c 3 1 c 0 0 a
2 79 40 c0011 5 10 203cc 77 78 32 0 11aa aa aa aa aa aa aa aa
2 80 40 70008 0 1 400 0 0 x6
2 81 40 70011 3 35 f00e 79 80
2 82 41 120012 5 1 c 0 0 b
2 83 41 d000d 3 1 c 0 0 a
2 84 41 d0012 5 11 203cc 82 83 1 0 1102
2 85 41 70009 0 1 400 0 0 w10
2 86 41 70012 3 35 f00e 84 85
2 87 42 130013 5 1 c 0 0 b
2 88 42 d000d 3 1 c 0 0 a
2 89 42 d0013 5 12 203cc 87 88 1 0 1102
2 90 42 70009 0 1 400 0 0 w11
2 91 42 70013 3 35 f00e 89 90
2 92 43 120012 5 1 c 0 0 b
2 93 43 d000d 3 1 c 0 0 a
2 94 43 d0012 5 13 203cc 92 93 1 0 1102
2 95 43 70009 0 1 400 0 0 w12
2 96 43 70012 3 35 f00e 94 95
2 97 44 120012 5 1 c 0 0 b
2 98 44 d000d 3 1 c 0 0 a
2 99 44 d0012 5 14 203cc 97 98 1 0 1102
2 100 44 70009 0 1 400 0 0 w13
2 101 44 70012 3 35 f00e 99 100
2 102 45 120012 5 1 c 0 0 b
2 103 45 d000d 3 1 c 0 0 a
2 104 45 d0012 5 15 203cc 102 103 1 0 1102
2 105 45 70009 0 1 400 0 0 w14
2 106 45 70012 3 35 f00e 104 105
2 107 46 130013 5 1 c 0 0 b
2 108 46 d000d 3 1 c 0 0 a
2 109 46 d0013 5 16 203cc 107 108 1 0 1102
2 110 46 70009 0 1 400 0 0 w15
2 111 46 70013 3 35 f00e 109 110
2 112 47 120012 5 1 c 0 0 b
2 113 47 d000d 3 1 c 0 0 a
2 114 47 d0012 5 17 203cc 112 113 1 0 1102
2 115 47 70009 0 1 400 0 0 w16
2 116 47 70012 3 35 f00e 114 115
2 117 48 120012 5 1 c 0 0 b
2 118 48 d000d 3 1 c 0 0 a
2 119 48 d0012 5 18 203cc 117 118 1 0 1102
2 120 48 70009 0 1 400 0 0 w17
2 121 48 70012 3 35 f00e 119 120
2 122 49 150015 8 1 c 0 0 c
2 123 49 110011 5 1 c 0 0 b
2 124 49 d0011 9 1a 203cc 122 123 1 0 1102
2 125 49 d000d 3 1 c 0 0 a
2 126 49 d0015 9 19 203cc 124 125 1 0 1102
2 127 49 70009 0 1 400 0 0 w18
2 128 49 70015 6 35 f00e 126 127
2 129 50 e000e 3 1 c 0 0 a
2 130 50 d000d 3 1b 2000c 129 0 1 0 1102
2 131 50 70009 0 1 400 0 0 w19
2 132 50 7000e 3 35 f00e 130 131
2 133 51 e000e 40 1 c 0 0 d
2 134 51 d000d 40 1c 2000c 133 0 1 0 1102
2 135 51 70009 0 1 400 0 0 w20
2 136 51 7000e 10 35 f00e 134 135
2 137 52 e000e 3 1 c 0 0 a
2 138 52 d000d 3 1d 2000c 137 0 1 0 1102
2 139 52 70009 0 1 400 0 0 w21
2 140 52 7000e 3 35 f00e 138 139
2 141 53 e000e 40 1 c 0 0 d
2 142 53 d000d 40 1e 2000c 141 0 1 0 1102
2 143 53 70009 0 1 400 0 0 w22
2 144 53 7000e 10 35 f00e 142 143
2 145 54 e000e 40 1 c 0 0 d
2 146 54 d000d 40 1f 2000c 145 0 1 0 1102
2 147 54 70009 0 1 400 0 0 w23
2 148 54 7000e 30 35 f00e 146 147
2 149 55 f000f 40 1 c 0 0 d
2 150 55 d000e 40 20 2000c 149 0 1 0 1102
2 151 55 70009 0 1 400 0 0 w24
2 152 55 7000f 11 35 f00e 150 151
2 153 56 f000f 40 1 c 0 0 d
2 154 56 d000e 40 21 2000c 153 0 1 0 1102
2 155 56 70009 0 1 400 0 0 w25
2 156 56 7000f 11 35 f00e 154 155
2 157 57 f000f 40 1 c 0 0 d
2 158 57 d000e 40 22 2000c 157 0 1 0 1102
2 159 57 70009 0 1 400 0 0 w26
2 160 57 7000f 30 35 f00e 158 159
2 161 58 f000f 41 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 162 58 d0010 41 23 c 0 161 d
2 163 58 70009 0 1 400 0 0 w27
2 164 58 70010 41 35 f00e 162 163
2 165 59 110011 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 166 59 f000f 41 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 167 59 d0012 41 24 20c 165 166 d
2 168 59 70008 0 1 400 0 0 y0
2 169 59 70012 41 35 f00e 167 168
2 170 60 100010 3 1 c 0 0 a
2 171 60 e000e 1 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 172 60 d0012 4 25 2030c 170 171 2 0 330a
2 173 60 70008 0 1 400 0 0 y1
2 174 60 70012 4 35 f00e 172 173
2 175 61 110011 5 1 c 0 0 b
2 176 61 e000e 3 1 c 0 0 a
2 177 61 e0011 5 31 203cc 175 176 2 0 330a
2 178 61 d0012 5 26 2000c 177 0 2 0 330a
2 179 61 70008 0 1 400 0 0 y2
2 180 61 70012 5 35 f00e 178 179
1 a 0 3 30008 1 0 1102
1 b 0 3 3000b 1 0 1102
1 c 0 3 3000e 1 0 1102
1 d 0 4 3000c 3 0 772a
1 w0 0 6 3000c 1 0 2
1 w1 0 7 3000c 1 0 1102
1 w2 0 7 30010 1 0 1102
1 w3 0 7 30014 1 0 1102
1 w4 0 7 30018 1 0 1102
1 w5 0 8 3000c 1 0 1102
1 w6 0 9 3000c 1 0 1102
1 w7 0 10 3000c 1 0 1102
1 w8 0 10 30010 1 0 1102
1 w9 0 10 30014 1 0 1102
1 w10 0 11 3000c 1 0 1102
1 w11 0 11 30011 1 0 1102
1 w12 0 11 30016 1 0 1102
1 w13 0 11 3001b 1 0 1102
1 w14 0 11 30020 1 0 1102
1 w15 0 11 30025 1 0 1102
1 w16 0 11 3002a 1 0 1102
1 w17 0 11 3002f 1 0 1102
1 w18 0 11 30034 1 0 1102
1 w19 0 11 30039 1 0 1102
1 w20 0 12 3000c 1 0 1102
1 w21 0 12 30011 1 0 1102
1 w22 0 12 30016 1 0 1102
1 w23 0 12 3001b 1 0 1102
1 w24 0 12 30020 1 0 1102
1 w25 0 12 30025 1 0 1102
1 w26 0 12 3002a 1 0 1102
1 w27 0 12 3002f 1 0 1102
1 x0 0 13 3000c 32 0 11aa aa aa aa aa aa aa aa
1 x1 0 14 3000c 32 0 11aa aa aa aa aa aa aa aa
1 x2 0 15 3000c 32 0 11aa aa aa aa aa aa aa aa
1 x3 0 16 3000c 32 0 33aa aa aa aa aa aa aa aa
1 x4 0 16 30010 32 0 ffaa ffaa ffaa ffaa ffaa ffaa ffaa ffaa
1 x5 0 16 30014 32 0 33aa aa aa aa aa aa aa aa
1 x6 0 16 30018 32 0 11aa aa aa aa aa aa aa aa
1 y0 0 17 3000c 2 0 330a
1 y1 0 18 3000c 2 0 330a
1 y2 0 19 3000c 2 0 330a
1 i 0 21 3000c 32 96 13aa aa aa aa aa aa aa aa
1 j 0 22 3000c 32 96 13aa aa aa aa aa aa aa aa
1 k 0 22 3000f 32 96 13aa aa aa aa aa aa aa aa
1 l 0 22 30012 32 96 7faa aa aa aa aa aa aa aa
4 3 3 3
4 6 6 6
4 11 11 11
4 16 16 16
4 21 21 21
4 26 26 26
4 31 31 31
4 36 36 36
4 41 41 41
4 46 46 46
4 51 51 51
4 56 56 56
4 61 61 61
4 66 66 66
4 71 71 71
4 76 76 76
4 81 81 81
4 86 86 86
4 91 91 91
4 96 96 96
4 101 101 101
4 106 106 106
4 111 111 111
4 116 116 116
4 121 121 121
4 128 128 128
4 132 132 132
4 136 136 136
4 140 140 140
4 144 144 144
4 148 148 148
4 152 152 152
4 156 156 156
4 160 160 160
4 164 164 164
4 169 169 169
4 174 174 174
4 180 180 180
*/

/* OUTPUT assign1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : assign1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    assign1.v                 38/    0/   38      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    assign1.v                 79/  185/  264       30%            79/  185/  264       30%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: assign1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      w0                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x0                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x1                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x2                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x3                        0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0003 ...
      x5                        0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0003 ...
      x6                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              assign1.v                          96/   0/  96      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    assign1.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT assign1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : assign1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    assign1.v                 38/    0/   38      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    assign1.v                 79/  185/  264       30%            79/  185/  264       30%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: assign1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      w0                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x0                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x1                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x2                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x3                        0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0003 ...
      x5                        0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0003 ...
      x6                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              assign1.v                          96/   0/  96      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    assign1.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT assign1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : assign1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         38/    0/   38      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         79/  185/  264       30%            79/  185/  264       30%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: assign1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      w0                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x0                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x1                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x2                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x3                        0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0003 ...
      x5                        0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0003 ...
      x6                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            96/   0/  96      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT assign1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : assign1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         38/    0/   38      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         79/  185/  264       30%            79/  185/  264       30%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: assign1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      w0                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x0                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x1                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x2                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...
      x3                        0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0003 ...
      x5                        0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0003 ...
      x6                        0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0001 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            96/   0/  96      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
