module main;

parameter STATE_IDLE = 2'b00,
          STATE_HEAD = 2'b01,
          STATE_DATA = 2'b10,
          STATE_TAIL = 2'b11;

reg        clk;
reg        reset;
reg        head;
reg        tail;
reg        valid;
reg [1:0]  state;
reg [1:0]  next_state;

always @(posedge clk) state <= reset ? STATE_IDLE : next_state;

(* covered_fsm, channel, is="state", os="next_state",
                         trans="STATE_HEAD->STATE_DATA",
                         trans="STATE_DATA->STATE_TAIL",
                         trans="STATE_DATA->STATE_DATA",
                         trans="STATE_TAIL->STATE_HEAD" *)
always @(state or head or valid or tail)
  begin
   case( state )
     STATE_IDLE:  next_state = (valid & head) ? STATE_HEAD : STATE_IDLE;
     STATE_HEAD:  next_state = (valid & tail) ? STATE_TAIL : STATE_DATA;
     STATE_DATA:  next_state = (valid & tail) ? STATE_TAIL : STATE_DATA;
     STATE_TAIL:  next_state = (valid & head) ? STATE_HEAD : STATE_IDLE;
   endcase
  end

initial begin
	$dumpfile( "fsm7.3.vcd" );
	$dumpvars( 0, main );
        reset = 1'b1;
	head  = 1'b0;
        tail  = 1'b0;
        valid = 1'b0;
	#20;
	reset = 1'b0;
	#20;
	@(posedge clk);
        head <= 1'b1;
	valid <= 1'b1;
	@(posedge clk);
        head <= 1'b0;
	tail <= 1'b1;
	@(posedge clk);
	tail  <= 1'b0;
	valid <= 1'b0;
	#20;
	$finish;
end

initial begin
	clk = 1'b0;
        forever #(2) clk = ~clk;
end

endmodule

/* HEADER
GROUPS fsm7.3 all iv vcd lxt
SIM    fsm7.3 all iv vcd  : iverilog fsm7.3.v; ./a.out                             : fsm7.3.vcd
SIM    fsm7.3 all iv lxt  : iverilog fsm7.3.v; ./a.out -lxt2; mv fsm7.3.vcd fsm7.3.lxt : fsm7.3.lxt
SCORE  fsm7.3.vcd     : -t main -vcd fsm7.3.vcd -o fsm7.3.cdd -v fsm7.3.v : fsm7.3.cdd
SCORE  fsm7.3.lxt     : -t main -lxt fsm7.3.lxt -o fsm7.3.cdd -v fsm7.3.v : fsm7.3.cdd
REPORT fsm7.3.cdd 1   : -d v -o fsm7.3.rptM fsm7.3.cdd                         : fsm7.3.rptM
REPORT fsm7.3.cdd 2   : -d v -w -o fsm7.3.rptWM fsm7.3.cdd                     : fsm7.3.rptWM
REPORT fsm7.3.cdd 3   : -d v -i -o fsm7.3.rptI fsm7.3.cdd                      : fsm7.3.rptI
REPORT fsm7.3.cdd 4   : -d v -w -i -o fsm7.3.rptWI fsm7.3.cdd                  : fsm7.3.rptWI
*/

/* OUTPUT fsm7.3.cdd
5 1 * 6 0 0 0 0
3 0 main main fsm7.3.v 1 61
2 1 16 34003d 5 1 c 0 0 next_state
2 2 16 270030 1 32 4 0 0 #STATE_IDLE
2 3 16 1f0030 7 1a 200cc 1 2 32 0 33aa aa aa aa aa aa aa aa
2 4 16 1f0023 2 1 c 0 0 reset
2 5 16 1f003d 7 19 201cc 3 4 2 0 330a
2 6 16 16001a 0 1 400 0 0 state
2 7 16 16003d 12 38 600e 5 6
2 8 16 110013 24 1 c 0 0 clk
2 9 16 9000f 0 2a 20000 0 0 2 0 a
2 10 16 90013 37 27 2100a 8 9 1 0 2
2 11 26 3d0046 1 32 4 0 0 #STATE_IDLE
2 12 26 300039 1 32 8 0 0 #STATE_HEAD
2 13 26 1f0039 3 1a 2010c 11 12 32 0 11aa aa aa aa aa aa aa aa
2 14 26 28002b 3 1 c 0 0 head
2 15 26 200024 3 1 c 0 0 valid
2 16 26 20002b 3 8 2024c 14 15 1 0 1102
2 17 26 1f0046 3 19 2024c 13 16 2 0 110a
2 18 26 12001b 0 1 400 0 0 next_state
2 19 26 120046 3 37 600e 17 18
2 20 27 3d0046 1 32 8 0 0 #STATE_DATA
2 21 27 300039 1 32 8 0 0 #STATE_TAIL
2 22 27 1f0039 1 1a 20208 20 21 32 0 aa aa aa aa aa aa aa aa
2 23 27 28002b 1 1 18 0 0 tail
2 24 27 200024 1 1 18 0 0 valid
2 25 27 20002b 1 8 20238 23 24 1 0 2
2 26 27 1f0046 1 19 20238 22 25 2 0 a
2 27 27 12001b 0 1 400 0 0 next_state
2 28 27 120046 1 37 602a 26 27
2 29 28 3d0046 0 32 10 0 0 #STATE_DATA
2 30 28 300039 0 32 10 0 0 #STATE_TAIL
2 31 28 1f0039 0 1a 20030 29 30 32 0 aa aa aa aa aa aa aa aa
2 32 28 28002b 0 1 10 0 0 tail
2 33 28 200024 0 1 10 0 0 valid
2 34 28 20002b 0 8 20030 32 33 1 0 2
2 35 28 1f0046 0 19 20030 31 34 2 0 a
2 36 28 12001b 0 1 400 0 0 next_state
2 37 28 120046 0 37 6022 35 36
2 38 29 3d0046 1 32 4 0 0 #STATE_IDLE
2 39 29 300039 1 32 8 0 0 #STATE_HEAD
2 40 29 1f0039 1 1a 20104 38 39 32 0 aa aa aa aa aa aa aa aa
2 41 29 28002b 1 1 4 0 0 head
2 42 29 200024 1 1 4 0 0 valid
2 43 29 20002b 1 8 20044 41 42 1 0 2
2 44 29 1f0046 1 19 20044 40 43 2 0 a
2 45 29 12001b 0 1 400 0 0 next_state
2 46 29 120046 1 37 6006 44 45
2 47 29 5000e 1 32 8 0 0 #STATE_TAIL
2 48 25 9000d d 1 e 0 0 state
2 49 29 0 2 2d 2420e 47 48 1 0 102
2 50 28 5000e 1 32 8 0 0 #STATE_DATA
2 51 28 0 2 2d 20206 50 48 1 0 2
2 52 27 5000e 1 32 8 0 0 #STATE_HEAD
2 53 27 0 3 2d 2020e 52 48 1 0 1102
2 54 26 5000e 1 32 4 0 0 #STATE_IDLE
2 55 26 0 6 2d 2014e 54 48 1 0 1102
2 56 23 230026 3 1 c 0 0 tail
2 57 23 230026 0 2a 20000 0 0 2 0 110a
2 58 23 230026 3 29 20008 56 57 1 0 2
2 59 23 1a001e 3 1 c 0 0 valid
2 60 23 1a001e 0 2a 20000 0 0 2 0 110a
2 61 23 1a001e 3 29 20008 59 60 1 0 2
2 62 23 120015 3 1 c 0 0 head
2 63 23 120015 0 2a 20000 0 0 2 0 110a
2 64 23 120015 3 29 20008 62 63 1 0 2
2 65 23 9000d 5 1 c 0 0 state
2 66 23 9000d 0 2a 20000 0 0 3 0 332a
2 67 23 9000d 5 29 20008 65 66 1 0 2
2 68 23 90015 6 2b 20008 64 67 1 0 2
2 69 23 9001e 6 2b 20008 61 68 1 0 2
2 70 23 90026 d 2b 2100a 58 69 1 0 2
2 71 57 7000a 1 0 20004 0 0 1 1 0
2 72 57 10003 0 1 400 0 0 clk
2 73 57 1000a 1 37 1006 71 72
2 74 58 1c001e 23 1 1c 0 0 clk
2 75 58 1b001b 23 1b 2002c 74 0 1 0 1102
2 76 58 150017 0 1 400 0 0 clk
2 77 58 15001e 23 37 602e 75 76
2 78 58 120012 1 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 79 58 120012 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 80 58 100013 47 2c 2000a 78 79 32 0 aa aa aa aa aa aa aa aa
2 81 0 0 5 1 f00e 0 0 next_state
2 82 0 0 5 1 f00e 0 0 state
1 #STATE_IDLE 0 0 0 32 0 0 0 0 0 0 0 0 0
1 #STATE_HEAD 0 0 0 32 0 1 0 0 0 0 0 0 0
1 #STATE_DATA 0 0 0 32 0 4 0 0 0 0 0 0 0
1 #STATE_TAIL 0 0 0 32 0 5 0 0 0 0 0 0 0
1 clk 0 8 3000b 1 16 1102
1 reset 0 9 3000b 1 0 1002
1 head 0 10 3000b 1 0 1102
1 tail 0 11 3000b 1 0 1102
1 valid 0 12 3000b 1 0 1102
1 state 0 13 3000b 2 0 330a
1 next_state 0 14 3000b 2 16 330a
4 82 82 82
4 81 81 81
4 7 10 10
4 10 7 0
4 46 70 70
4 49 46 70
4 37 70 70
4 51 37 49
4 28 70 70
4 53 28 51
4 19 70 70
4 55 19 53
4 70 55 0
4 77 80 80
4 80 77 0
4 73 80 80
6 82 81 1 02,08,08,01c0,60014001a00101,21,e1,8101
*/

/* OUTPUT fsm7.3.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm7.3.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.3.v                   8/    1/    9       89%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           28:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.3.v                   8/    1/    9       89%             9/    0/    9      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm7.3.v                           21/  16/  37       57%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.3.v                  3/   1/   4       75%            4/   4/   8       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          2'h2

        Missed State Transitions

          From State    To State  
          ==========    ==========
          2'h1       -> 2'h2      
          2'h2       -> 2'h3      
          2'h2       -> 2'h2      
          2'h3       -> 2'h1      



*/

/* OUTPUT fsm7.3.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm7.3.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.3.v                   8/    1/    9       89%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           28:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.3.v                   8/    1/    9       89%             9/    0/    9      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm7.3.v                           21/  16/  37       57%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.3.v                  3/   1/   4       75%            4/   4/   8       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          2'h2

        Missed State Transitions

          From State    To State  
          ==========    ==========
          2'h1       -> 2'h2      
          2'h2       -> 2'h3      
          2'h2       -> 2'h2      
          2'h3       -> 2'h1      



*/

/* OUTPUT fsm7.3.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm7.3.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          8/    1/    9       89%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           28:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          8/    1/    9       89%             9/    0/    9      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            21/  16/  37       57%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         3/   1/   4       75%            4/   4/   8       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          2'h2

        Missed State Transitions

          From State    To State  
          ==========    ==========
          2'h1       -> 2'h2      
          2'h2       -> 2'h3      
          2'h2       -> 2'h2      
          2'h3       -> 2'h1      



*/

/* OUTPUT fsm7.3.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm7.3.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          8/    1/    9       89%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           28:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          8/    1/    9       89%             9/    0/    9      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            21/  16/  37       57%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         3/   1/   4       75%            4/   4/   8       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          2'h2

        Missed State Transitions

          From State    To State  
          ==========    ==========
          2'h1       -> 2'h2      
          2'h2       -> 2'h3      
          2'h2       -> 2'h2      
          2'h3       -> 2'h1      



*/
