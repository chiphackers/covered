module main;

foo f( 1'b0 );

endmodule

//--------------------------

module foo (
  input wire a
);

endmodule
