module main;

wire        a;
reg         b, c;
reg  [27:3] d;
reg         e;

assign a = (b | c) &
                   ((d[27:16]==12'h0) &&
                    (d[12:3] != 10'h000) &&
                    (d[12:3] != 10'h001) &&
                    (d[12:3] != 10'h002) &&
                    (d[12:3] != 10'h003) &&
                    (d[12:3] != 10'h004) &&
                    (d[12:3] != 10'h005) &&
                    (d[12:3] != 10'h006) &&
                    (d[12:3] != 10'h007) &&
                    (d[12:3] != 10'h008) &&
                    (d[12:3] != 10'h009) &&
                    (d[12:3] != 10'h00A) &&
                    (d[12:3] != 10'h00B) &&
                    (d[12:3] != 10'h00C) &&
                    (d[12:3] != 10'h00D) &&
                    (d[12:3] != 10'h00E) &&
                    (d[12:3] != 10'h00F) &&
                    (d[12:3] != 10'h010) &&
                    (d[12:3] != 10'h011) &&
                    (d[12:3] != 10'h012) &&
                    (d[12:3] != 10'h013) &&
                    (d[12:3] != 10'h014) &&
                    (d[12:3] != 10'h015) &&
                    (d[12:3] != 10'h016) &&
                    (d[12:3] != 10'h017) &&
                    (d[12:3] != 10'h018) &&
                    (d[12:3] != 10'h019) &&
                    (d[12:3] != 10'h01A) &&
                    (d[12:3] != 10'h01B) &&
                    (d[12:3] != 10'h01C) &&
                    (d[12:3] != 10'h01D) &&
                    (d[12:3] != 10'h01E) &&
                    (d[12:3] != 10'h01F) &&
                    (d[12:3] != 10'h020) &&
                    (d[12:3] != 10'h021) &&
                    (d[12:3] != 10'h022) &&
                    (d[12:3] != 10'h023) &&
                    (d[12:3] != 10'h024) &&
                    (d[12:3] != 10'h025) &&
                    (d[12:3] != 10'h026) &&
                    (d[12:3] != 10'h027) &&
                    (d[12:3] != 10'h028) &&
                    (d[12:3] != 10'h029) &&
                    (d[12:3] != 10'h02A) &&
                    (d[12:3] != 10'h02B) &&
                    (d[12:3] != 10'h02C) &&
                    (d[12:3] != 10'h02D) &&
                    (d[12:3] != 10'h02E) &&
                    (d[12:3] != 10'h02F) &&
                    (d[12:3] != 10'h030) &&
                    (d[12:3] != 10'h031) &&
                    (d[12:3] != 10'h032) &&
                    (d[12:3] != 10'h033) &&
                    (d[12:3] != 10'h034) &&
                    (d[12:3] != 10'h035) &&
                    (d[12:3] != 10'h036) &&
                    (d[12:3] != 10'h037) &&
                    (d[12:3] != 10'h038) &&
                    (d[12:3] != 10'h039) &&
                    (d[12:3] != 10'h03A) &&
                    (d[12:3] != 10'h03B) &&
                    (d[12:3] != 10'h03C) &&
                    (d[12:3] != 10'h03D) &&
                    (d[12:3] != 10'h03E) &&
                    (d[12:3] != 10'h03F) &&
                    (d[12:3] != 10'h040) &&
                    (d[12:3] != 10'h041) &&
                    (d[12:3] != 10'h042) &&
                    (d[12:3] != 10'h043) &&
                    (d[12:3] != 10'h044) &&
                    (d[12:3] != 10'h045) &&
                    (d[12:3] != 10'h046) &&
                    (d[12:3] != 10'h047) &&
                    (d[12:3] != 10'h048) &&
                    (d[12:3] != 10'h049) &&
                    (d[12:3] != 10'h04A) &&
                    (d[12:3] != 10'h04B) &&
                    (d[12:3] != 10'h04C) &&
                    (d[12:3] != 10'h04D) &&
                    (d[12:3] != 10'h04E) &&
                    (d[12:3] != 10'h04F) &&
                    (d[12:3] != 10'h050) &&
                    (d[12:3] != 10'h051) &&
                    (d[12:3] != 10'h052) &&
                    (d[12:3] != 10'h053) &&
                    (d[12:3] != 10'h054)) |
                   e &
                   ((d[27:16]==12'h0) &&
                    (d[12:3] != 10'h000) &&
                    (d[12:3] != 10'h001) &&
                    (d[12:3] != 10'h002) &&
                    (d[12:3] != 10'h003) &&
                    (d[12:3] != 10'h004) &&
                    (d[12:3] != 10'h005) &&
                    (d[12:3] != 10'h006) &&
                    (d[12:3] != 10'h007) &&
                    (d[12:3] != 10'h008) &&
                    (d[12:3] != 10'h009) &&
                    (d[12:3] != 10'h00A) &&
                    (d[12:3] != 10'h00B) &&
                    (d[12:3] != 10'h00C) &&
                    (d[12:3] != 10'h00D) &&
                    (d[12:3] != 10'h00E) &&
                    (d[12:3] != 10'h00F) &&
                    (d[12:3] != 10'h010) &&
                    (d[12:3] != 10'h011) &&
                    (d[12:3] != 10'h012) &&
                    (d[12:3] != 10'h013) &&
                    (d[12:3] != 10'h014) &&
                    (d[12:3] != 10'h015) &&
                    (d[12:3] != 10'h016) &&
                    (d[12:3] != 10'h017) &&
                    (d[12:3] != 10'h018) &&
                    (d[12:3] != 10'h019) &&
                    (d[12:3] != 10'h01A) &&
                    (d[12:3] != 10'h01B) &&
                    (d[12:3] != 10'h01C) &&
                    (d[12:3] != 10'h01D) &&
                    (d[12:3] != 10'h01E) &&
                    (d[12:3] != 10'h01F) &&
                    (d[12:3] != 10'h020) &&
                    (d[12:3] != 10'h021) &&
                    (d[12:3] != 10'h022) &&
                    (d[12:3] != 10'h023) &&
                    (d[12:3] != 10'h024) &&
                    (d[12:3] != 10'h025) &&
                    (d[12:3] != 10'h026) &&
                    (d[12:3] != 10'h027) &&
                    (d[12:3] != 10'h028) &&
                    (d[12:3] != 10'h029) &&
                    (d[12:3] != 10'h02A) &&
                    (d[12:3] != 10'h02B) &&
                    (d[12:3] != 10'h02C) &&
                    (d[12:3] != 10'h02D) &&
                    (d[12:3] != 10'h02E) &&
                    (d[12:3] != 10'h02F) &&
                    (d[12:3] != 10'h030) &&
                    (d[12:3] != 10'h031) &&
                    (d[12:3] != 10'h032) &&
                    (d[12:3] != 10'h033) &&
                    (d[12:3] != 10'h034) &&
                    (d[12:3] != 10'h035) &&
                    (d[12:3] != 10'h036) &&
                    (d[12:3] != 10'h037) &&
                    (d[12:3] != 10'h038) &&
                    (d[12:3] != 10'h039) &&
                    (d[12:3] != 10'h03A) &&
                    (d[12:3] != 10'h03B) &&
                    (d[12:3] != 10'h03C) &&
                    (d[12:3] != 10'h03D) &&
                    (d[12:3] != 10'h03E) &&
                    (d[12:3] != 10'h03F) &&
                    (d[12:3] != 10'h040) &&
                    (d[12:3] != 10'h041) &&
                    (d[12:3] != 10'h042) &&
                    (d[12:3] != 10'h043) &&
                    (d[12:3] != 10'h044) &&
                    (d[12:3] != 10'h045) &&
                    (d[12:3] != 10'h046) &&
                    (d[12:3] != 10'h047) &&
                    (d[12:3] != 10'h048) &&
                    (d[12:3] != 10'h049) &&
                    (d[12:3] != 10'h04A) &&
                    (d[12:3] != 10'h04B)) ;

initial begin
	$dumpfile( "long_exp1.vcd" );
	$dumpvars( 0, main );
	b = 1'b0;
	c = 1'b0;
	d = 25'h0000000;
	e = 1'b0;
	#5;
	$finish;
end

endmodule

/* HEADER
GROUPS long_exp1 all iv vcs vcd lxt
SIM    long_exp1 all iv vcd  : iverilog long_exp1.v; ./a.out                             : long_exp1.vcd
SIM    long_exp1 all iv lxt  : iverilog long_exp1.v; ./a.out -lxt2; mv long_exp1.vcd long_exp1.lxt : long_exp1.lxt
SIM    long_exp1 all vcs vcd : vcs long_exp1.v; ./simv                                   : long_exp1.vcd
SCORE  long_exp1.vcd     : -t main -vcd long_exp1.vcd -o long_exp1.cdd -v long_exp1.v : long_exp1.cdd
SCORE  long_exp1.lxt     : -t main -lxt long_exp1.lxt -o long_exp1.cdd -v long_exp1.v : long_exp1.cdd
REPORT long_exp1.cdd 1   : -d v -o long_exp1.rptM long_exp1.cdd                         : long_exp1.rptM
REPORT long_exp1.cdd 2   : -d v -w -o long_exp1.rptWM long_exp1.cdd                     : long_exp1.rptWM
REPORT long_exp1.cdd 3   : -d v -i -o long_exp1.rptI long_exp1.cdd                      : long_exp1.rptI
REPORT long_exp1.cdd 4   : -d v -w -i -o long_exp1.rptWI long_exp1.cdd                  : long_exp1.rptWI
*/

/* OUTPUT long_exp1.cdd
5 1 * 6 0 0 0 0
3 0 main main long_exp1.v 1 185
2 1 172 200026 1 0 20008 0 0 10 3 45 10 0
2 2 172 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 3 172 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 4 172 15001b 2 24 204 2 3 d
2 5 172 150026 2 15 20088 1 4 1 0 2
2 6 171 200026 1 0 20008 0 0 10 3 44 10 0
2 7 171 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 8 171 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 9 171 15001b 2 24 204 7 8 d
2 10 171 150026 2 15 20088 6 9 1 0 2
2 11 170 200026 1 0 20008 0 0 10 3 41 10 0
2 12 170 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 13 170 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 14 170 15001b 2 24 204 12 13 d
2 15 170 150026 2 15 20088 11 14 1 0 2
2 16 169 200026 1 0 20008 0 0 10 3 40 10 0
2 17 169 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 18 169 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 19 169 15001b 2 24 204 17 18 d
2 20 169 150026 2 15 20088 16 19 1 0 2
2 21 168 200026 1 0 20008 0 0 10 3 15 10 0
2 22 168 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 23 168 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 24 168 15001b 2 24 204 22 23 d
2 25 168 150026 2 15 20088 21 24 1 0 2
2 26 167 200026 1 0 20008 0 0 10 3 14 10 0
2 27 167 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 28 167 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 29 167 15001b 2 24 204 27 28 d
2 30 167 150026 2 15 20088 26 29 1 0 2
2 31 166 200026 1 0 20008 0 0 10 3 11 10 0
2 32 166 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 33 166 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 34 166 15001b 2 24 204 32 33 d
2 35 166 150026 2 15 20088 31 34 1 0 2
2 36 165 200026 1 0 20008 0 0 10 3 10 10 0
2 37 165 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 38 165 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 39 165 15001b 2 24 204 37 38 d
2 40 165 150026 2 15 20088 36 39 1 0 2
2 41 164 200026 1 0 20008 0 0 10 3 5 10 0
2 42 164 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 43 164 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 44 164 15001b 2 24 204 42 43 d
2 45 164 150026 2 15 20088 41 44 1 0 2
2 46 163 200026 1 0 20008 0 0 10 3 4 10 0
2 47 163 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 48 163 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 49 163 15001b 2 24 204 47 48 d
2 50 163 150026 2 15 20088 46 49 1 0 2
2 51 162 200026 1 0 20008 0 0 10 3 1 10 0
2 52 162 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 53 162 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 54 162 15001b 2 24 204 52 53 d
2 55 162 150026 2 15 20088 51 54 1 0 2
2 56 161 200026 1 0 20008 0 0 10 3 0 10 0
2 57 161 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 58 161 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 59 161 15001b 2 24 204 57 58 d
2 60 161 150026 2 15 20088 56 59 1 0 2
2 61 160 200026 1 0 20008 0 0 10 3 55 5 0
2 62 160 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 63 160 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 64 160 15001b 2 24 204 62 63 d
2 65 160 150026 2 15 20088 61 64 1 0 2
2 66 159 200026 1 0 20008 0 0 10 3 54 5 0
2 67 159 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 68 159 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 69 159 15001b 2 24 204 67 68 d
2 70 159 150026 2 15 20088 66 69 1 0 2
2 71 158 200026 1 0 20008 0 0 10 3 51 5 0
2 72 158 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 73 158 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 74 158 15001b 2 24 204 72 73 d
2 75 158 150026 2 15 20088 71 74 1 0 2
2 76 157 200026 1 0 20008 0 0 10 3 50 5 0
2 77 157 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 78 157 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 79 157 15001b 2 24 204 77 78 d
2 80 157 150026 2 15 20088 76 79 1 0 2
2 81 156 200026 1 0 20008 0 0 10 3 45 5 0
2 82 156 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 83 156 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 84 156 15001b 2 24 204 82 83 d
2 85 156 150026 2 15 20088 81 84 1 0 2
2 86 155 200026 1 0 20008 0 0 10 3 44 5 0
2 87 155 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 88 155 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 89 155 15001b 2 24 204 87 88 d
2 90 155 150026 2 15 20088 86 89 1 0 2
2 91 154 200026 1 0 20008 0 0 10 3 41 5 0
2 92 154 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 93 154 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 94 154 15001b 2 24 204 92 93 d
2 95 154 150026 2 15 20088 91 94 1 0 2
2 96 153 200026 1 0 20008 0 0 10 3 40 5 0
2 97 153 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 98 153 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 99 153 15001b 2 24 204 97 98 d
2 100 153 150026 2 15 20088 96 99 1 0 2
2 101 152 200026 1 0 20008 0 0 10 3 15 5 0
2 102 152 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 103 152 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 104 152 15001b 2 24 204 102 103 d
2 105 152 150026 2 15 20088 101 104 1 0 2
2 106 151 200026 1 0 20008 0 0 10 3 14 5 0
2 107 151 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 108 151 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 109 151 15001b 2 24 204 107 108 d
2 110 151 150026 2 15 20088 106 109 1 0 2
2 111 150 200026 1 0 20008 0 0 10 3 11 5 0
2 112 150 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 113 150 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 114 150 15001b 2 24 204 112 113 d
2 115 150 150026 2 15 20088 111 114 1 0 2
2 116 149 200026 1 0 20008 0 0 10 3 10 5 0
2 117 149 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 118 149 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 119 149 15001b 2 24 204 117 118 d
2 120 149 150026 2 15 20088 116 119 1 0 2
2 121 148 200026 1 0 20008 0 0 10 3 5 5 0
2 122 148 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 123 148 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 124 148 15001b 2 24 204 122 123 d
2 125 148 150026 2 15 20088 121 124 1 0 2
2 126 147 200026 1 0 20008 0 0 10 3 4 5 0
2 127 147 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 128 147 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 129 147 15001b 2 24 204 127 128 d
2 130 147 150026 2 15 20088 126 129 1 0 2
2 131 146 200026 1 0 20008 0 0 10 3 1 5 0
2 132 146 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 133 146 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 134 146 15001b 2 24 204 132 133 d
2 135 146 150026 2 15 20088 131 134 1 0 2
2 136 145 200026 1 0 20008 0 0 10 3 0 5 0
2 137 145 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 138 145 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 139 145 15001b 2 24 204 137 138 d
2 140 145 150026 2 15 20088 136 139 1 0 2
2 141 144 200026 1 0 20008 0 0 10 3 55 4 0
2 142 144 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 143 144 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 144 144 15001b 2 24 204 142 143 d
2 145 144 150026 2 15 20088 141 144 1 0 2
2 146 143 200026 1 0 20008 0 0 10 3 54 4 0
2 147 143 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 148 143 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 149 143 15001b 2 24 204 147 148 d
2 150 143 150026 2 15 20088 146 149 1 0 2
2 151 142 200026 1 0 20008 0 0 10 3 51 4 0
2 152 142 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 153 142 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 154 142 15001b 2 24 204 152 153 d
2 155 142 150026 2 15 20088 151 154 1 0 2
2 156 141 200026 1 0 20008 0 0 10 3 50 4 0
2 157 141 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 158 141 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 159 141 15001b 2 24 204 157 158 d
2 160 141 150026 2 15 20088 156 159 1 0 2
2 161 140 200026 1 0 20008 0 0 10 3 45 4 0
2 162 140 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 163 140 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 164 140 15001b 2 24 204 162 163 d
2 165 140 150026 2 15 20088 161 164 1 0 2
2 166 139 200026 1 0 20008 0 0 10 3 44 4 0
2 167 139 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 168 139 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 169 139 15001b 2 24 204 167 168 d
2 170 139 150026 2 15 20088 166 169 1 0 2
2 171 138 200026 1 0 20008 0 0 10 3 41 4 0
2 172 138 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 173 138 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 174 138 15001b 2 24 204 172 173 d
2 175 138 150026 2 15 20088 171 174 1 0 2
2 176 137 200026 1 0 20008 0 0 10 3 40 4 0
2 177 137 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 178 137 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 179 137 15001b 2 24 204 177 178 d
2 180 137 150026 2 15 20088 176 179 1 0 2
2 181 136 200026 1 0 20008 0 0 10 3 15 4 0
2 182 136 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 183 136 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 184 136 15001b 2 24 204 182 183 d
2 185 136 150026 2 15 20088 181 184 1 0 2
2 186 135 200026 1 0 20008 0 0 10 3 14 4 0
2 187 135 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 188 135 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 189 135 15001b 2 24 204 187 188 d
2 190 135 150026 2 15 20088 186 189 1 0 2
2 191 134 200026 1 0 20008 0 0 10 3 11 4 0
2 192 134 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 193 134 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 194 134 15001b 2 24 204 192 193 d
2 195 134 150026 2 15 20088 191 194 1 0 2
2 196 133 200026 1 0 20008 0 0 10 3 10 4 0
2 197 133 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 198 133 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 199 133 15001b 2 24 204 197 198 d
2 200 133 150026 2 15 20088 196 199 1 0 2
2 201 132 200026 1 0 20008 0 0 10 3 5 4 0
2 202 132 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 203 132 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 204 132 15001b 2 24 204 202 203 d
2 205 132 150026 2 15 20088 201 204 1 0 2
2 206 131 200026 1 0 20008 0 0 10 3 4 4 0
2 207 131 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 208 131 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 209 131 15001b 2 24 204 207 208 d
2 210 131 150026 2 15 20088 206 209 1 0 2
2 211 130 200026 1 0 20008 0 0 10 3 1 4 0
2 212 130 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 213 130 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 214 130 15001b 2 24 204 212 213 d
2 215 130 150026 2 15 20088 211 214 1 0 2
2 216 129 200026 1 0 20008 0 0 10 3 0 4 0
2 217 129 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 218 129 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 219 129 15001b 2 24 204 217 218 d
2 220 129 150026 2 15 20088 216 219 1 0 2
2 221 128 200026 1 0 20008 0 0 10 3 55 1 0
2 222 128 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 223 128 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 224 128 15001b 2 24 204 222 223 d
2 225 128 150026 2 15 20088 221 224 1 0 2
2 226 127 200026 1 0 20008 0 0 10 3 54 1 0
2 227 127 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 228 127 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 229 127 15001b 2 24 204 227 228 d
2 230 127 150026 2 15 20088 226 229 1 0 2
2 231 126 200026 1 0 20008 0 0 10 3 51 1 0
2 232 126 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 233 126 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 234 126 15001b 2 24 204 232 233 d
2 235 126 150026 2 15 20088 231 234 1 0 2
2 236 125 200026 1 0 20008 0 0 10 3 50 1 0
2 237 125 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 238 125 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 239 125 15001b 2 24 204 237 238 d
2 240 125 150026 2 15 20088 236 239 1 0 2
2 241 124 200026 1 0 20008 0 0 10 3 45 1 0
2 242 124 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 243 124 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 244 124 15001b 2 24 204 242 243 d
2 245 124 150026 2 15 20088 241 244 1 0 2
2 246 123 200026 1 0 20008 0 0 10 3 44 1 0
2 247 123 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 248 123 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 249 123 15001b 2 24 204 247 248 d
2 250 123 150026 2 15 20088 246 249 1 0 2
2 251 122 200026 1 0 20008 0 0 10 3 41 1 0
2 252 122 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 253 122 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 254 122 15001b 2 24 204 252 253 d
2 255 122 150026 2 15 20088 251 254 1 0 2
2 256 121 200026 1 0 20008 0 0 10 3 40 1 0
2 257 121 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 258 121 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 259 121 15001b 2 24 204 257 258 d
2 260 121 150026 2 15 20088 256 259 1 0 2
2 261 120 200026 1 0 20008 0 0 10 3 15 1 0
2 262 120 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 263 120 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 264 120 15001b 2 24 204 262 263 d
2 265 120 150026 2 15 20088 261 264 1 0 2
2 266 119 200026 1 0 20008 0 0 10 3 14 1 0
2 267 119 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 268 119 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 269 119 15001b 2 24 204 267 268 d
2 270 119 150026 2 15 20088 266 269 1 0 2
2 271 118 200026 1 0 20008 0 0 10 3 11 1 0
2 272 118 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 273 118 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 274 118 15001b 2 24 204 272 273 d
2 275 118 150026 2 15 20088 271 274 1 0 2
2 276 117 200026 1 0 20008 0 0 10 3 10 1 0
2 277 117 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 278 117 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 279 117 15001b 2 24 204 277 278 d
2 280 117 150026 2 15 20088 276 279 1 0 2
2 281 116 200026 1 0 20008 0 0 10 3 5 1 0
2 282 116 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 283 116 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 284 116 15001b 2 24 204 282 283 d
2 285 116 150026 2 15 20088 281 284 1 0 2
2 286 115 200026 1 0 20008 0 0 10 3 4 1 0
2 287 115 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 288 115 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 289 115 15001b 2 24 204 287 288 d
2 290 115 150026 2 15 20088 286 289 1 0 2
2 291 114 200026 1 0 20008 0 0 10 3 1 1 0
2 292 114 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 293 114 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 294 114 15001b 2 24 204 292 293 d
2 295 114 150026 2 15 20088 291 294 1 0 2
2 296 113 200026 1 0 20008 0 0 10 3 0 1 0
2 297 113 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 298 113 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 299 113 15001b 2 24 204 297 298 d
2 300 113 150026 2 15 20088 296 299 1 0 2
2 301 112 200026 1 0 20008 0 0 10 3 55 0 0
2 302 112 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 303 112 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 304 112 15001b 2 24 204 302 303 d
2 305 112 150026 2 15 20088 301 304 1 0 2
2 306 111 200026 1 0 20008 0 0 10 3 54 0 0
2 307 111 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 308 111 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 309 111 15001b 2 24 204 307 308 d
2 310 111 150026 2 15 20088 306 309 1 0 2
2 311 110 200026 1 0 20008 0 0 10 3 51 0 0
2 312 110 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 313 110 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 314 110 15001b 2 24 204 312 313 d
2 315 110 150026 2 15 20088 311 314 1 0 2
2 316 109 200026 1 0 20008 0 0 10 3 50 0 0
2 317 109 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 318 109 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 319 109 15001b 2 24 204 317 318 d
2 320 109 150026 2 15 20088 316 319 1 0 2
2 321 108 200026 1 0 20008 0 0 10 3 45 0 0
2 322 108 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 323 108 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 324 108 15001b 2 24 204 322 323 d
2 325 108 150026 2 15 20088 321 324 1 0 2
2 326 107 200026 1 0 20008 0 0 10 3 44 0 0
2 327 107 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 328 107 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 329 107 15001b 2 24 204 327 328 d
2 330 107 150026 2 15 20088 326 329 1 0 2
2 331 106 200026 1 0 20008 0 0 10 3 41 0 0
2 332 106 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 333 106 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 334 106 15001b 2 24 204 332 333 d
2 335 106 150026 2 15 20088 331 334 1 0 2
2 336 105 200026 1 0 20008 0 0 10 3 40 0 0
2 337 105 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 338 105 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 339 105 15001b 2 24 204 337 338 d
2 340 105 150026 2 15 20088 336 339 1 0 2
2 341 104 200026 1 0 20008 0 0 10 3 15 0 0
2 342 104 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 343 104 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 344 104 15001b 2 24 204 342 343 d
2 345 104 150026 2 15 20088 341 344 1 0 2
2 346 103 200026 1 0 20008 0 0 10 3 14 0 0
2 347 103 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 348 103 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 349 103 15001b 2 24 204 347 348 d
2 350 103 150026 2 15 20088 346 349 1 0 2
2 351 102 200026 1 0 20008 0 0 10 3 11 0 0
2 352 102 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 353 102 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 354 102 15001b 2 24 204 352 353 d
2 355 102 150026 2 15 20088 351 354 1 0 2
2 356 101 200026 1 0 20008 0 0 10 3 10 0 0
2 357 101 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 358 101 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 359 101 15001b 2 24 204 357 358 d
2 360 101 150026 2 15 20088 356 359 1 0 2
2 361 100 200026 1 0 20008 0 0 10 3 5 0 0
2 362 100 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 363 100 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 364 100 15001b 2 24 204 362 363 d
2 365 100 150026 2 15 20088 361 364 1 0 2
2 366 99 200026 1 0 20008 0 0 10 3 4 0 0
2 367 99 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 368 99 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 369 99 15001b 2 24 204 367 368 d
2 370 99 150026 2 15 20088 366 369 1 0 2
2 371 98 200026 1 0 20008 0 0 10 3 1 0 0
2 372 98 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 373 98 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 374 98 15001b 2 24 204 372 373 d
2 375 98 150026 2 15 20088 371 374 1 0 2
2 376 97 200026 1 0 20004 0 0 10 3 0 0 0
2 377 97 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 378 97 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 379 97 15001b 2 24 204 377 378 d
2 380 97 150026 2 15 20044 376 379 1 0 2
2 381 96 1f0023 1 0 20004 0 0 12 3 0 0 0
2 382 96 1a001b 1 0 20008 0 0 32 64 0 1 0 0 0 0 0 0
2 383 96 170018 2 0 20008 0 0 32 64 45 1 0 0 0 0 0 0
2 384 96 15001c 2 24 204 382 383 d
2 385 96 150023 2 11 20048 381 384 1 0 2
2 386 96 140027 2 18 20104 380 385 1 0 2
2 387 96 140027 2 18 20084 375 386 1 0 2
2 388 96 140027 2 18 20084 370 387 1 0 2
2 389 96 140027 2 18 20084 365 388 1 0 2
2 390 96 140027 2 18 20084 360 389 1 0 2
2 391 96 140027 2 18 20084 355 390 1 0 2
2 392 96 140027 2 18 20084 350 391 1 0 2
2 393 96 140027 2 18 20084 345 392 1 0 2
2 394 96 140027 2 18 20084 340 393 1 0 2
2 395 96 140027 2 18 20084 335 394 1 0 2
2 396 96 140027 2 18 20084 330 395 1 0 2
2 397 96 140027 2 18 20084 325 396 1 0 2
2 398 96 140027 2 18 20084 320 397 1 0 2
2 399 96 140027 2 18 20084 315 398 1 0 2
2 400 96 140027 2 18 20084 310 399 1 0 2
2 401 96 140027 2 18 20084 305 400 1 0 2
2 402 96 140027 2 18 20084 300 401 1 0 2
2 403 96 140027 2 18 20084 295 402 1 0 2
2 404 96 140027 2 18 20084 290 403 1 0 2
2 405 96 140027 2 18 20084 285 404 1 0 2
2 406 96 140027 2 18 20084 280 405 1 0 2
2 407 96 140027 2 18 20084 275 406 1 0 2
2 408 96 140027 2 18 20084 270 407 1 0 2
2 409 96 140027 2 18 20084 265 408 1 0 2
2 410 96 140027 2 18 20084 260 409 1 0 2
2 411 96 140027 2 18 20084 255 410 1 0 2
2 412 96 140027 2 18 20084 250 411 1 0 2
2 413 96 140027 2 18 20084 245 412 1 0 2
2 414 96 140027 2 18 20084 240 413 1 0 2
2 415 96 140027 2 18 20084 235 414 1 0 2
2 416 96 140027 2 18 20084 230 415 1 0 2
2 417 96 140027 2 18 20084 225 416 1 0 2
2 418 96 140027 2 18 20084 220 417 1 0 2
2 419 96 140027 2 18 20084 215 418 1 0 2
2 420 96 140027 2 18 20084 210 419 1 0 2
2 421 96 140027 2 18 20084 205 420 1 0 2
2 422 96 140027 2 18 20084 200 421 1 0 2
2 423 96 140027 2 18 20084 195 422 1 0 2
2 424 96 140027 2 18 20084 190 423 1 0 2
2 425 96 140027 2 18 20084 185 424 1 0 2
2 426 96 140027 2 18 20084 180 425 1 0 2
2 427 96 140027 2 18 20084 175 426 1 0 2
2 428 96 140027 2 18 20084 170 427 1 0 2
2 429 96 140027 2 18 20084 165 428 1 0 2
2 430 96 140027 2 18 20084 160 429 1 0 2
2 431 96 140027 2 18 20084 155 430 1 0 2
2 432 96 140027 2 18 20084 150 431 1 0 2
2 433 96 140027 2 18 20084 145 432 1 0 2
2 434 96 140027 2 18 20084 140 433 1 0 2
2 435 96 140027 2 18 20084 135 434 1 0 2
2 436 96 140027 2 18 20084 130 435 1 0 2
2 437 96 140027 2 18 20084 125 436 1 0 2
2 438 96 140027 2 18 20084 120 437 1 0 2
2 439 96 140027 2 18 20084 115 438 1 0 2
2 440 96 140027 2 18 20084 110 439 1 0 2
2 441 96 140027 2 18 20084 105 440 1 0 2
2 442 96 140027 2 18 20084 100 441 1 0 2
2 443 96 140027 2 18 20084 95 442 1 0 2
2 444 96 140027 2 18 20084 90 443 1 0 2
2 445 96 140027 2 18 20084 85 444 1 0 2
2 446 96 140027 2 18 20084 80 445 1 0 2
2 447 96 140027 2 18 20084 75 446 1 0 2
2 448 96 140027 2 18 20084 70 447 1 0 2
2 449 96 140027 2 18 20084 65 448 1 0 2
2 450 96 140027 2 18 20084 60 449 1 0 2
2 451 96 140027 2 18 20084 55 450 1 0 2
2 452 96 140027 2 18 20084 50 451 1 0 2
2 453 96 140027 2 18 20084 45 452 1 0 2
2 454 96 140027 2 18 20084 40 453 1 0 2
2 455 96 140027 2 18 20084 35 454 1 0 2
2 456 96 140027 2 18 20084 30 455 1 0 2
2 457 96 140027 2 18 20084 25 456 1 0 2
2 458 96 140027 2 18 20084 20 457 1 0 2
2 459 96 140027 2 18 20084 15 458 1 0 2
2 460 96 140027 2 18 20084 10 459 1 0 2
2 461 96 140027 2 18 20084 5 460 1 0 2
2 462 95 130013 1 1 4 0 0 e
2 463 95 130028 2 8 20044 461 462 1 0 2
2 464 94 200026 1 0 20008 0 0 10 3 10 11 0
2 465 94 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 466 94 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 467 94 15001b 2 24 204 465 466 d
2 468 94 150026 2 15 20088 464 467 1 0 2
2 469 93 200026 1 0 20008 0 0 10 3 5 11 0
2 470 93 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 471 93 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 472 93 15001b 2 24 204 470 471 d
2 473 93 150026 2 15 20088 469 472 1 0 2
2 474 92 200026 1 0 20008 0 0 10 3 4 11 0
2 475 92 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 476 92 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 477 92 15001b 2 24 204 475 476 d
2 478 92 150026 2 15 20088 474 477 1 0 2
2 479 91 200026 1 0 20008 0 0 10 3 1 11 0
2 480 91 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 481 91 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 482 91 15001b 2 24 204 480 481 d
2 483 91 150026 2 15 20088 479 482 1 0 2
2 484 90 200026 1 0 20008 0 0 10 3 0 11 0
2 485 90 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 486 90 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 487 90 15001b 2 24 204 485 486 d
2 488 90 150026 2 15 20088 484 487 1 0 2
2 489 89 200026 1 0 20008 0 0 10 3 55 10 0
2 490 89 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 491 89 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 492 89 15001b 2 24 204 490 491 d
2 493 89 150026 2 15 20088 489 492 1 0 2
2 494 88 200026 1 0 20008 0 0 10 3 54 10 0
2 495 88 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 496 88 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 497 88 15001b 2 24 204 495 496 d
2 498 88 150026 2 15 20088 494 497 1 0 2
2 499 87 200026 1 0 20008 0 0 10 3 51 10 0
2 500 87 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 501 87 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 502 87 15001b 2 24 204 500 501 d
2 503 87 150026 2 15 20088 499 502 1 0 2
2 504 86 200026 1 0 20008 0 0 10 3 50 10 0
2 505 86 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 506 86 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 507 86 15001b 2 24 204 505 506 d
2 508 86 150026 2 15 20088 504 507 1 0 2
2 509 85 200026 1 0 20008 0 0 10 3 45 10 0
2 510 85 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 511 85 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 512 85 15001b 2 24 204 510 511 d
2 513 85 150026 2 15 20088 509 512 1 0 2
2 514 84 200026 1 0 20008 0 0 10 3 44 10 0
2 515 84 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 516 84 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 517 84 15001b 2 24 204 515 516 d
2 518 84 150026 2 15 20088 514 517 1 0 2
2 519 83 200026 1 0 20008 0 0 10 3 41 10 0
2 520 83 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 521 83 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 522 83 15001b 2 24 204 520 521 d
2 523 83 150026 2 15 20088 519 522 1 0 2
2 524 82 200026 1 0 20008 0 0 10 3 40 10 0
2 525 82 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 526 82 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 527 82 15001b 2 24 204 525 526 d
2 528 82 150026 2 15 20088 524 527 1 0 2
2 529 81 200026 1 0 20008 0 0 10 3 15 10 0
2 530 81 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 531 81 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 532 81 15001b 2 24 204 530 531 d
2 533 81 150026 2 15 20088 529 532 1 0 2
2 534 80 200026 1 0 20008 0 0 10 3 14 10 0
2 535 80 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 536 80 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 537 80 15001b 2 24 204 535 536 d
2 538 80 150026 2 15 20088 534 537 1 0 2
2 539 79 200026 1 0 20008 0 0 10 3 11 10 0
2 540 79 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 541 79 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 542 79 15001b 2 24 204 540 541 d
2 543 79 150026 2 15 20088 539 542 1 0 2
2 544 78 200026 1 0 20008 0 0 10 3 10 10 0
2 545 78 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 546 78 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 547 78 15001b 2 24 204 545 546 d
2 548 78 150026 2 15 20088 544 547 1 0 2
2 549 77 200026 1 0 20008 0 0 10 3 5 10 0
2 550 77 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 551 77 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 552 77 15001b 2 24 204 550 551 d
2 553 77 150026 2 15 20088 549 552 1 0 2
2 554 76 200026 1 0 20008 0 0 10 3 4 10 0
2 555 76 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 556 76 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 557 76 15001b 2 24 204 555 556 d
2 558 76 150026 2 15 20088 554 557 1 0 2
2 559 75 200026 1 0 20008 0 0 10 3 1 10 0
2 560 75 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 561 75 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 562 75 15001b 2 24 204 560 561 d
2 563 75 150026 2 15 20088 559 562 1 0 2
2 564 74 200026 1 0 20008 0 0 10 3 0 10 0
2 565 74 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 566 74 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 567 74 15001b 2 24 204 565 566 d
2 568 74 150026 2 15 20088 564 567 1 0 2
2 569 73 200026 1 0 20008 0 0 10 3 55 5 0
2 570 73 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 571 73 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 572 73 15001b 2 24 204 570 571 d
2 573 73 150026 2 15 20088 569 572 1 0 2
2 574 72 200026 1 0 20008 0 0 10 3 54 5 0
2 575 72 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 576 72 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 577 72 15001b 2 24 204 575 576 d
2 578 72 150026 2 15 20088 574 577 1 0 2
2 579 71 200026 1 0 20008 0 0 10 3 51 5 0
2 580 71 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 581 71 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 582 71 15001b 2 24 204 580 581 d
2 583 71 150026 2 15 20088 579 582 1 0 2
2 584 70 200026 1 0 20008 0 0 10 3 50 5 0
2 585 70 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 586 70 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 587 70 15001b 2 24 204 585 586 d
2 588 70 150026 2 15 20088 584 587 1 0 2
2 589 69 200026 1 0 20008 0 0 10 3 45 5 0
2 590 69 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 591 69 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 592 69 15001b 2 24 204 590 591 d
2 593 69 150026 2 15 20088 589 592 1 0 2
2 594 68 200026 1 0 20008 0 0 10 3 44 5 0
2 595 68 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 596 68 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 597 68 15001b 2 24 204 595 596 d
2 598 68 150026 2 15 20088 594 597 1 0 2
2 599 67 200026 1 0 20008 0 0 10 3 41 5 0
2 600 67 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 601 67 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 602 67 15001b 2 24 204 600 601 d
2 603 67 150026 2 15 20088 599 602 1 0 2
2 604 66 200026 1 0 20008 0 0 10 3 40 5 0
2 605 66 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 606 66 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 607 66 15001b 2 24 204 605 606 d
2 608 66 150026 2 15 20088 604 607 1 0 2
2 609 65 200026 1 0 20008 0 0 10 3 15 5 0
2 610 65 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 611 65 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 612 65 15001b 2 24 204 610 611 d
2 613 65 150026 2 15 20088 609 612 1 0 2
2 614 64 200026 1 0 20008 0 0 10 3 14 5 0
2 615 64 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 616 64 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 617 64 15001b 2 24 204 615 616 d
2 618 64 150026 2 15 20088 614 617 1 0 2
2 619 63 200026 1 0 20008 0 0 10 3 11 5 0
2 620 63 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 621 63 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 622 63 15001b 2 24 204 620 621 d
2 623 63 150026 2 15 20088 619 622 1 0 2
2 624 62 200026 1 0 20008 0 0 10 3 10 5 0
2 625 62 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 626 62 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 627 62 15001b 2 24 204 625 626 d
2 628 62 150026 2 15 20088 624 627 1 0 2
2 629 61 200026 1 0 20008 0 0 10 3 5 5 0
2 630 61 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 631 61 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 632 61 15001b 2 24 204 630 631 d
2 633 61 150026 2 15 20088 629 632 1 0 2
2 634 60 200026 1 0 20008 0 0 10 3 4 5 0
2 635 60 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 636 60 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 637 60 15001b 2 24 204 635 636 d
2 638 60 150026 2 15 20088 634 637 1 0 2
2 639 59 200026 1 0 20008 0 0 10 3 1 5 0
2 640 59 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 641 59 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 642 59 15001b 2 24 204 640 641 d
2 643 59 150026 2 15 20088 639 642 1 0 2
2 644 58 200026 1 0 20008 0 0 10 3 0 5 0
2 645 58 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 646 58 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 647 58 15001b 2 24 204 645 646 d
2 648 58 150026 2 15 20088 644 647 1 0 2
2 649 57 200026 1 0 20008 0 0 10 3 55 4 0
2 650 57 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 651 57 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 652 57 15001b 2 24 204 650 651 d
2 653 57 150026 2 15 20088 649 652 1 0 2
2 654 56 200026 1 0 20008 0 0 10 3 54 4 0
2 655 56 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 656 56 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 657 56 15001b 2 24 204 655 656 d
2 658 56 150026 2 15 20088 654 657 1 0 2
2 659 55 200026 1 0 20008 0 0 10 3 51 4 0
2 660 55 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 661 55 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 662 55 15001b 2 24 204 660 661 d
2 663 55 150026 2 15 20088 659 662 1 0 2
2 664 54 200026 1 0 20008 0 0 10 3 50 4 0
2 665 54 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 666 54 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 667 54 15001b 2 24 204 665 666 d
2 668 54 150026 2 15 20088 664 667 1 0 2
2 669 53 200026 1 0 20008 0 0 10 3 45 4 0
2 670 53 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 671 53 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 672 53 15001b 2 24 204 670 671 d
2 673 53 150026 2 15 20088 669 672 1 0 2
2 674 52 200026 1 0 20008 0 0 10 3 44 4 0
2 675 52 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 676 52 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 677 52 15001b 2 24 204 675 676 d
2 678 52 150026 2 15 20088 674 677 1 0 2
2 679 51 200026 1 0 20008 0 0 10 3 41 4 0
2 680 51 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 681 51 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 682 51 15001b 2 24 204 680 681 d
2 683 51 150026 2 15 20088 679 682 1 0 2
2 684 50 200026 1 0 20008 0 0 10 3 40 4 0
2 685 50 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 686 50 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 687 50 15001b 2 24 204 685 686 d
2 688 50 150026 2 15 20088 684 687 1 0 2
2 689 49 200026 1 0 20008 0 0 10 3 15 4 0
2 690 49 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 691 49 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 692 49 15001b 2 24 204 690 691 d
2 693 49 150026 2 15 20088 689 692 1 0 2
2 694 48 200026 1 0 20008 0 0 10 3 14 4 0
2 695 48 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 696 48 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 697 48 15001b 2 24 204 695 696 d
2 698 48 150026 2 15 20088 694 697 1 0 2
2 699 47 200026 1 0 20008 0 0 10 3 11 4 0
2 700 47 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 701 47 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 702 47 15001b 2 24 204 700 701 d
2 703 47 150026 2 15 20088 699 702 1 0 2
2 704 46 200026 1 0 20008 0 0 10 3 10 4 0
2 705 46 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 706 46 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 707 46 15001b 2 24 204 705 706 d
2 708 46 150026 2 15 20088 704 707 1 0 2
2 709 45 200026 1 0 20008 0 0 10 3 5 4 0
2 710 45 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 711 45 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 712 45 15001b 2 24 204 710 711 d
2 713 45 150026 2 15 20088 709 712 1 0 2
2 714 44 200026 1 0 20008 0 0 10 3 4 4 0
2 715 44 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 716 44 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 717 44 15001b 2 24 204 715 716 d
2 718 44 150026 2 15 20088 714 717 1 0 2
2 719 43 200026 1 0 20008 0 0 10 3 1 4 0
2 720 43 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 721 43 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 722 43 15001b 2 24 204 720 721 d
2 723 43 150026 2 15 20088 719 722 1 0 2
2 724 42 200026 1 0 20008 0 0 10 3 0 4 0
2 725 42 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 726 42 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 727 42 15001b 2 24 204 725 726 d
2 728 42 150026 2 15 20088 724 727 1 0 2
2 729 41 200026 1 0 20008 0 0 10 3 55 1 0
2 730 41 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 731 41 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 732 41 15001b 2 24 204 730 731 d
2 733 41 150026 2 15 20088 729 732 1 0 2
2 734 40 200026 1 0 20008 0 0 10 3 54 1 0
2 735 40 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 736 40 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 737 40 15001b 2 24 204 735 736 d
2 738 40 150026 2 15 20088 734 737 1 0 2
2 739 39 200026 1 0 20008 0 0 10 3 51 1 0
2 740 39 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 741 39 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 742 39 15001b 2 24 204 740 741 d
2 743 39 150026 2 15 20088 739 742 1 0 2
2 744 38 200026 1 0 20008 0 0 10 3 50 1 0
2 745 38 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 746 38 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 747 38 15001b 2 24 204 745 746 d
2 748 38 150026 2 15 20088 744 747 1 0 2
2 749 37 200026 1 0 20008 0 0 10 3 45 1 0
2 750 37 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 751 37 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 752 37 15001b 2 24 204 750 751 d
2 753 37 150026 2 15 20088 749 752 1 0 2
2 754 36 200026 1 0 20008 0 0 10 3 44 1 0
2 755 36 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 756 36 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 757 36 15001b 2 24 204 755 756 d
2 758 36 150026 2 15 20088 754 757 1 0 2
2 759 35 200026 1 0 20008 0 0 10 3 41 1 0
2 760 35 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 761 35 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 762 35 15001b 2 24 204 760 761 d
2 763 35 150026 2 15 20088 759 762 1 0 2
2 764 34 200026 1 0 20008 0 0 10 3 40 1 0
2 765 34 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 766 34 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 767 34 15001b 2 24 204 765 766 d
2 768 34 150026 2 15 20088 764 767 1 0 2
2 769 33 200026 1 0 20008 0 0 10 3 15 1 0
2 770 33 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 771 33 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 772 33 15001b 2 24 204 770 771 d
2 773 33 150026 2 15 20088 769 772 1 0 2
2 774 32 200026 1 0 20008 0 0 10 3 14 1 0
2 775 32 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 776 32 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 777 32 15001b 2 24 204 775 776 d
2 778 32 150026 2 15 20088 774 777 1 0 2
2 779 31 200026 1 0 20008 0 0 10 3 11 1 0
2 780 31 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 781 31 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 782 31 15001b 2 24 204 780 781 d
2 783 31 150026 2 15 20088 779 782 1 0 2
2 784 30 200026 1 0 20008 0 0 10 3 10 1 0
2 785 30 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 786 30 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 787 30 15001b 2 24 204 785 786 d
2 788 30 150026 2 15 20088 784 787 1 0 2
2 789 29 200026 1 0 20008 0 0 10 3 5 1 0
2 790 29 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 791 29 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 792 29 15001b 2 24 204 790 791 d
2 793 29 150026 2 15 20088 789 792 1 0 2
2 794 28 200026 1 0 20008 0 0 10 3 4 1 0
2 795 28 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 796 28 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 797 28 15001b 2 24 204 795 796 d
2 798 28 150026 2 15 20088 794 797 1 0 2
2 799 27 200026 1 0 20008 0 0 10 3 1 1 0
2 800 27 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 801 27 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 802 27 15001b 2 24 204 800 801 d
2 803 27 150026 2 15 20088 799 802 1 0 2
2 804 26 200026 1 0 20008 0 0 10 3 0 1 0
2 805 26 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 806 26 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 807 26 15001b 2 24 204 805 806 d
2 808 26 150026 2 15 20088 804 807 1 0 2
2 809 25 200026 1 0 20008 0 0 10 3 55 0 0
2 810 25 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 811 25 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 812 25 15001b 2 24 204 810 811 d
2 813 25 150026 2 15 20088 809 812 1 0 2
2 814 24 200026 1 0 20008 0 0 10 3 54 0 0
2 815 24 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 816 24 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 817 24 15001b 2 24 204 815 816 d
2 818 24 150026 2 15 20088 814 817 1 0 2
2 819 23 200026 1 0 20008 0 0 10 3 51 0 0
2 820 23 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 821 23 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 822 23 15001b 2 24 204 820 821 d
2 823 23 150026 2 15 20088 819 822 1 0 2
2 824 22 200026 1 0 20008 0 0 10 3 50 0 0
2 825 22 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 826 22 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 827 22 15001b 2 24 204 825 826 d
2 828 22 150026 2 15 20088 824 827 1 0 2
2 829 21 200026 1 0 20008 0 0 10 3 45 0 0
2 830 21 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 831 21 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 832 21 15001b 2 24 204 830 831 d
2 833 21 150026 2 15 20088 829 832 1 0 2
2 834 20 200026 1 0 20008 0 0 10 3 44 0 0
2 835 20 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 836 20 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 837 20 15001b 2 24 204 835 836 d
2 838 20 150026 2 15 20088 834 837 1 0 2
2 839 19 200026 1 0 20008 0 0 10 3 41 0 0
2 840 19 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 841 19 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 842 19 15001b 2 24 204 840 841 d
2 843 19 150026 2 15 20088 839 842 1 0 2
2 844 18 200026 1 0 20008 0 0 10 3 40 0 0
2 845 18 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 846 18 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 847 18 15001b 2 24 204 845 846 d
2 848 18 150026 2 15 20088 844 847 1 0 2
2 849 17 200026 1 0 20008 0 0 10 3 15 0 0
2 850 17 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 851 17 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 852 17 15001b 2 24 204 850 851 d
2 853 17 150026 2 15 20088 849 852 1 0 2
2 854 16 200026 1 0 20008 0 0 10 3 14 0 0
2 855 16 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 856 16 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 857 16 15001b 2 24 204 855 856 d
2 858 16 150026 2 15 20088 854 857 1 0 2
2 859 15 200026 1 0 20008 0 0 10 3 11 0 0
2 860 15 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 861 15 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 862 15 15001b 2 24 204 860 861 d
2 863 15 150026 2 15 20088 859 862 1 0 2
2 864 14 200026 1 0 20008 0 0 10 3 10 0 0
2 865 14 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 866 14 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 867 14 15001b 2 24 204 865 866 d
2 868 14 150026 2 15 20088 864 867 1 0 2
2 869 13 200026 1 0 20008 0 0 10 3 5 0 0
2 870 13 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 871 13 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 872 13 15001b 2 24 204 870 871 d
2 873 13 150026 2 15 20088 869 872 1 0 2
2 874 12 200026 1 0 20008 0 0 10 3 4 0 0
2 875 12 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 876 12 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 877 12 15001b 2 24 204 875 876 d
2 878 12 150026 2 15 20088 874 877 1 0 2
2 879 11 200026 1 0 20008 0 0 10 3 1 0 0
2 880 11 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 881 11 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 882 11 15001b 2 24 204 880 881 d
2 883 11 150026 2 15 20088 879 882 1 0 2
2 884 10 200026 1 0 20004 0 0 10 3 0 0 0
2 885 10 1a001a 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 886 10 170018 2 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 887 10 15001b 2 24 204 885 886 d
2 888 10 150026 2 15 20044 884 887 1 0 2
2 889 9 1f0023 1 0 20004 0 0 12 3 0 0 0
2 890 9 1a001b 1 0 20008 0 0 32 64 0 1 0 0 0 0 0 0
2 891 9 170018 2 0 20008 0 0 32 64 45 1 0 0 0 0 0 0
2 892 9 15001c 2 24 204 890 891 d
2 893 9 150023 2 11 20048 889 892 1 0 2
2 894 9 140027 2 18 20104 888 893 1 0 2
2 895 9 140027 2 18 20084 883 894 1 0 2
2 896 9 140027 2 18 20084 878 895 1 0 2
2 897 9 140027 2 18 20084 873 896 1 0 2
2 898 9 140027 2 18 20084 868 897 1 0 2
2 899 9 140027 2 18 20084 863 898 1 0 2
2 900 9 140027 2 18 20084 858 899 1 0 2
2 901 9 140027 2 18 20084 853 900 1 0 2
2 902 9 140027 2 18 20084 848 901 1 0 2
2 903 9 140027 2 18 20084 843 902 1 0 2
2 904 9 140027 2 18 20084 838 903 1 0 2
2 905 9 140027 2 18 20084 833 904 1 0 2
2 906 9 140027 2 18 20084 828 905 1 0 2
2 907 9 140027 2 18 20084 823 906 1 0 2
2 908 9 140027 2 18 20084 818 907 1 0 2
2 909 9 140027 2 18 20084 813 908 1 0 2
2 910 9 140027 2 18 20084 808 909 1 0 2
2 911 9 140027 2 18 20084 803 910 1 0 2
2 912 9 140027 2 18 20084 798 911 1 0 2
2 913 9 140027 2 18 20084 793 912 1 0 2
2 914 9 140027 2 18 20084 788 913 1 0 2
2 915 9 140027 2 18 20084 783 914 1 0 2
2 916 9 140027 2 18 20084 778 915 1 0 2
2 917 9 140027 2 18 20084 773 916 1 0 2
2 918 9 140027 2 18 20084 768 917 1 0 2
2 919 9 140027 2 18 20084 763 918 1 0 2
2 920 9 140027 2 18 20084 758 919 1 0 2
2 921 9 140027 2 18 20084 753 920 1 0 2
2 922 9 140027 2 18 20084 748 921 1 0 2
2 923 9 140027 2 18 20084 743 922 1 0 2
2 924 9 140027 2 18 20084 738 923 1 0 2
2 925 9 140027 2 18 20084 733 924 1 0 2
2 926 9 140027 2 18 20084 728 925 1 0 2
2 927 9 140027 2 18 20084 723 926 1 0 2
2 928 9 140027 2 18 20084 718 927 1 0 2
2 929 9 140027 2 18 20084 713 928 1 0 2
2 930 9 140027 2 18 20084 708 929 1 0 2
2 931 9 140027 2 18 20084 703 930 1 0 2
2 932 9 140027 2 18 20084 698 931 1 0 2
2 933 9 140027 2 18 20084 693 932 1 0 2
2 934 9 140027 2 18 20084 688 933 1 0 2
2 935 9 140027 2 18 20084 683 934 1 0 2
2 936 9 140027 2 18 20084 678 935 1 0 2
2 937 9 140027 2 18 20084 673 936 1 0 2
2 938 9 140027 2 18 20084 668 937 1 0 2
2 939 9 140027 2 18 20084 663 938 1 0 2
2 940 9 140027 2 18 20084 658 939 1 0 2
2 941 9 140027 2 18 20084 653 940 1 0 2
2 942 9 140027 2 18 20084 648 941 1 0 2
2 943 9 140027 2 18 20084 643 942 1 0 2
2 944 9 140027 2 18 20084 638 943 1 0 2
2 945 9 140027 2 18 20084 633 944 1 0 2
2 946 9 140027 2 18 20084 628 945 1 0 2
2 947 9 140027 2 18 20084 623 946 1 0 2
2 948 9 140027 2 18 20084 618 947 1 0 2
2 949 9 140027 2 18 20084 613 948 1 0 2
2 950 9 140027 2 18 20084 608 949 1 0 2
2 951 9 140027 2 18 20084 603 950 1 0 2
2 952 9 140027 2 18 20084 598 951 1 0 2
2 953 9 140027 2 18 20084 593 952 1 0 2
2 954 9 140027 2 18 20084 588 953 1 0 2
2 955 9 140027 2 18 20084 583 954 1 0 2
2 956 9 140027 2 18 20084 578 955 1 0 2
2 957 9 140027 2 18 20084 573 956 1 0 2
2 958 9 140027 2 18 20084 568 957 1 0 2
2 959 9 140027 2 18 20084 563 958 1 0 2
2 960 9 140027 2 18 20084 558 959 1 0 2
2 961 9 140027 2 18 20084 553 960 1 0 2
2 962 9 140027 2 18 20084 548 961 1 0 2
2 963 9 140027 2 18 20084 543 962 1 0 2
2 964 9 140027 2 18 20084 538 963 1 0 2
2 965 9 140027 2 18 20084 533 964 1 0 2
2 966 9 140027 2 18 20084 528 965 1 0 2
2 967 9 140027 2 18 20084 523 966 1 0 2
2 968 9 140027 2 18 20084 518 967 1 0 2
2 969 9 140027 2 18 20084 513 968 1 0 2
2 970 9 140027 2 18 20084 508 969 1 0 2
2 971 9 140027 2 18 20084 503 970 1 0 2
2 972 9 140027 2 18 20084 498 971 1 0 2
2 973 9 140027 2 18 20084 493 972 1 0 2
2 974 9 140027 2 18 20084 488 973 1 0 2
2 975 9 140027 2 18 20084 483 974 1 0 2
2 976 9 140027 2 18 20084 478 975 1 0 2
2 977 9 140027 2 18 20084 473 976 1 0 2
2 978 9 140027 2 18 20084 468 977 1 0 2
2 979 8 100010 1 1 4 0 0 c
2 980 8 c000c 1 1 4 0 0 b
2 981 8 c0010 1 9 20044 979 980 1 0 2
2 982 8 b0028 2 8 20044 978 981 1 0 2
2 983 8 b0028 2 9 20044 463 982 1 0 2
2 984 8 70007 0 1 400 0 0 a
2 985 8 70028 2 35 f006 983 984
1 a 0 3 3000c 1 0 2
1 b 0 4 3000c 1 0 2
1 c 0 4 3000f 1 0 2
1 d 3 5 3000c 25 0 aa aa aa aa aa aa 2
1 e 0 6 3000c 1 0 2
4 985 985 985
*/

/* OUTPUT long_exp1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : long_exp1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp1.v                1/    0/    1      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp1.v                0/   29/   29        0%             0/   29/   29        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 25'h000_0000
      ......................... 1->0: 25'h000_0000 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              long_exp1.v                       169/ 338/ 507       33%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              8:    assign  a  = ((( b  |  c ) & 
                                   |----1----|   
                                  |------89-------
                                 |------169-------
                    ((d[27:16] == 12'h0) && 
                     |--------2--------|    
                    |----------88------------
                    -----------89------------
                    -----------169-----------
                    (d[12:3] != 10'h0) && 
                    |-------3--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h1) && 
                    |-------4--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h2) && 
                    |-------5--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h3) && 
                    |-------6--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h4) && 
                    |-------7--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h5) && 
                    |-------8--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h6) && 
                    |-------9--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h7) && 
                    |-------10-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h8) && 
                    |-------11-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h9) && 
                    |-------12-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hA) && 
                    |-------13-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hB) && 
                    |-------14-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hC) && 
                    |-------15-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hD) && 
                    |-------16-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hE) && 
                    |-------17-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hF) && 
                    |-------18-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h10) && 
                    |-------19--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h11) && 
                    |-------20--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h12) && 
                    |-------21--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h13) && 
                    |-------22--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h14) && 
                    |-------23--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h15) && 
                    |-------24--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h16) && 
                    |-------25--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h17) && 
                    |-------26--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h18) && 
                    |-------27--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h19) && 
                    |-------28--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1A) && 
                    |-------29--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1B) && 
                    |-------30--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1C) && 
                    |-------31--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1D) && 
                    |-------32--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1E) && 
                    |-------33--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1F) && 
                    |-------34--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h20) && 
                    |-------35--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h21) && 
                    |-------36--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h22) && 
                    |-------37--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h23) && 
                    |-------38--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h24) && 
                    |-------39--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h25) && 
                    |-------40--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h26) && 
                    |-------41--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h27) && 
                    |-------42--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h28) && 
                    |-------43--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h29) && 
                    |-------44--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2A) && 
                    |-------45--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2B) && 
                    |-------46--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2C) && 
                    |-------47--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2D) && 
                    |-------48--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2E) && 
                    |-------49--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2F) && 
                    |-------50--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h30) && 
                    |-------51--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h31) && 
                    |-------52--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h32) && 
                    |-------53--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h33) && 
                    |-------54--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h34) && 
                    |-------55--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h35) && 
                    |-------56--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h36) && 
                    |-------57--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h37) && 
                    |-------58--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h38) && 
                    |-------59--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h39) && 
                    |-------60--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3A) && 
                    |-------61--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3B) && 
                    |-------62--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3C) && 
                    |-------63--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3D) && 
                    |-------64--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3E) && 
                    |-------65--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3F) && 
                    |-------66--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h40) && 
                    |-------67--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h41) && 
                    |-------68--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h42) && 
                    |-------69--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h43) && 
                    |-------70--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h44) && 
                    |-------71--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h45) && 
                    |-------72--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h46) && 
                    |-------73--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h47) && 
                    |-------74--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h48) && 
                    |-------75--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h49) && 
                    |-------76--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4A) && 
                    |-------77--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4B) && 
                    |-------78--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4C) && 
                    |-------79--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4D) && 
                    |-------80--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4E) && 
                    |-------81--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4F) && 
                    |-------82--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h50) && 
                    |-------83--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h51) && 
                    |-------84--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h52) && 
                    |-------85--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h53) && 
                    |-------86--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h54))) | 
                    |-------87--------|     
                    ---------88--------|    
                    ---------89---------|   
                    -----------169-----------
                    ( e  & 
                    |-168---
                    --169---
                    ((d[27:16] == 12'h0) && 
                     |-------90--------|    
                    |----------167-----------
                    -----------168-----------
                    -----------169-----------
                    (d[12:3] != 10'h0) && 
                    |-------91-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h1) && 
                    |-------92-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h2) && 
                    |-------93-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h3) && 
                    |-------94-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h4) && 
                    |-------95-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h5) && 
                    |-------96-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h6) && 
                    |-------97-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h7) && 
                    |-------98-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h8) && 
                    |-------99-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h9) && 
                    |------100-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hA) && 
                    |------101-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hB) && 
                    |------102-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hC) && 
                    |------103-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hD) && 
                    |------104-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hE) && 
                    |------105-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hF) && 
                    |------106-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h10) && 
                    |-------107-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h11) && 
                    |-------108-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h12) && 
                    |-------109-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h13) && 
                    |-------110-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h14) && 
                    |-------111-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h15) && 
                    |-------112-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h16) && 
                    |-------113-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h17) && 
                    |-------114-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h18) && 
                    |-------115-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h19) && 
                    |-------116-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1A) && 
                    |-------117-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1B) && 
                    |-------118-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1C) && 
                    |-------119-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1D) && 
                    |-------120-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1E) && 
                    |-------121-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1F) && 
                    |-------122-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h20) && 
                    |-------123-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h21) && 
                    |-------124-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h22) && 
                    |-------125-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h23) && 
                    |-------126-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h24) && 
                    |-------127-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h25) && 
                    |-------128-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h26) && 
                    |-------129-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h27) && 
                    |-------130-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h28) && 
                    |-------131-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h29) && 
                    |-------132-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2A) && 
                    |-------133-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2B) && 
                    |-------134-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2C) && 
                    |-------135-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2D) && 
                    |-------136-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2E) && 
                    |-------137-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2F) && 
                    |-------138-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h30) && 
                    |-------139-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h31) && 
                    |-------140-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h32) && 
                    |-------141-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h33) && 
                    |-------142-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h34) && 
                    |-------143-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h35) && 
                    |-------144-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h36) && 
                    |-------145-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h37) && 
                    |-------146-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h38) && 
                    |-------147-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h39) && 
                    |-------148-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3A) && 
                    |-------149-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3B) && 
                    |-------150-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3C) && 
                    |-------151-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3D) && 
                    |-------152-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3E) && 
                    |-------153-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3F) && 
                    |-------154-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h40) && 
                    |-------155-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h41) && 
                    |-------156-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h42) && 
                    |-------157-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h43) && 
                    |-------158-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h44) && 
                    |-------159-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h45) && 
                    |-------160-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h46) && 
                    |-------161-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h47) && 
                    |-------162-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h48) && 
                    |-------163-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h49) && 
                    |-------164-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h4A) && 
                    |-------165-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h4B))))
                    |-------166-------|   
                    --------167--------|  
                    ---------168--------| 
                    ---------169---------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 3   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
             *

        Expression 4   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 5   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 6   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 7   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 8   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 9   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 10   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 11   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 12   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 13   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 14   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 15   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 16   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 17   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 18   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 19   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 20   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 21   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 22   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 23   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 24   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 25   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 26   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 27   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 28   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 29   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 30   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 31   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 32   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 33   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 34   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 35   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 36   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 37   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 38   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 39   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 40   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 41   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 42   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 43   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 44   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 45   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 46   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 47   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 48   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 49   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 50   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 51   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 52   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 53   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 54   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 55   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 56   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 57   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 58   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 59   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 60   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 61   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 62   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 63   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 64   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 65   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 66   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 67   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 68   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 69   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 70   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 71   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 72   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 73   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 74   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 75   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 76   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 77   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 78   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 79   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 80   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 81   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 82   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 83   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 84   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 85   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 86   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 87   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 88   (1/87)
        ^^^^^^^^^^^^^ - &&
         2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 | 16 | 17 | 18 | 19 | 20 | 21 | 22 | 23 | 24 |
        =0=|=0=|=0=|=0=|=0=|=0=|=0=|=0=|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *       *   *   *   *   *   *   *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         25 | 26 | 27 | 28 | 29 | 30 | 31 | 32 | 33 | 34 | 35 | 36 | 37 | 38 | 39 | 40 | 41 | 42 | 43 | 44 | 45 | 46 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         47 | 48 | 49 | 50 | 51 | 52 | 53 | 54 | 55 | 56 | 57 | 58 | 59 | 60 | 61 | 62 | 63 | 64 | 65 | 66 | 67 | 68 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         69 | 70 | 71 | 72 | 73 | 74 | 75 | 76 | 77 | 78 | 79 | 80 | 81 | 82 | 83 | 84 | 85 | 86 | 87 | All
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|==1==
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *     *  

        Expression 89   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 90   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 91   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
             *

        Expression 92   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 93   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 94   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 95   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 96   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 97   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 98   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 99   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 100   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 101   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 102   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 103   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 104   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 105   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 106   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 107   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 108   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 109   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 110   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 111   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 112   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 113   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 114   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 115   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 116   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 117   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 118   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 119   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 120   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 121   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 122   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 123   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 124   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 125   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 126   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 127   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 128   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 129   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 130   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 131   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 132   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 133   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 134   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 135   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 136   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 137   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 138   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 139   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 140   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 141   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 142   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 143   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 144   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 145   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 146   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 147   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 148   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 149   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 150   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 151   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 152   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 153   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 154   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 155   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 156   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 157   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 158   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 159   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 160   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 161   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 162   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 163   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 164   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 165   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 166   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 167   (1/78)
        ^^^^^^^^^^^^^ - &&
         90 | 91 | 92 | 93 | 94 | 95 | 96 | 97 | 98 | 99 | 100 | 101 | 102 | 103 | 104 | 105 | 106 | 107 | 108 | 109 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *         *    *    *    *    *    *    *    *    *     *     *     *     *     *     *     *     *     *    

         110 | 111 | 112 | 113 | 114 | 115 | 116 | 117 | 118 | 119 | 120 | 121 | 122 | 123 | 124 | 125 | 126 | 127 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         128 | 129 | 130 | 131 | 132 | 133 | 134 | 135 | 136 | 137 | 138 | 139 | 140 | 141 | 142 | 143 | 144 | 145 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         146 | 147 | 148 | 149 | 150 | 151 | 152 | 153 | 154 | 155 | 156 | 157 | 158 | 159 | 160 | 161 | 162 | 163 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         164 | 165 | 166 | All
        =0===|=0===|=0===|==1==
         *     *     *      *  

        Expression 168   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 169   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp1.v               0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT long_exp1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : long_exp1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp1.v                1/    0/    1      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp1.v                0/   29/   29        0%             0/   29/   29        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 25'h000_0000
      ......................... 1->0: 25'h000_0000 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              long_exp1.v                       169/ 338/ 507       33%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              8:    assign  a  = ((( b  |  c ) & 
                                   |----1----|   
                                  |------89-------
                                 |------169-------
                    ((d[27:16] == 12'h0) && (d[12:3] != 10'h0) && (d[12:3] != 10'h1) && (d[12:3] != 10'h2) && 
                     |--------2--------|    |-------3--------|    |-------4--------|    |-------5--------|    
                    |-------------------------------------------88---------------------------------------------
                    --------------------------------------------89---------------------------------------------
                    --------------------------------------------169--------------------------------------------
                    (d[12:3] != 10'h3) && (d[12:3] != 10'h4) && (d[12:3] != 10'h5) && (d[12:3] != 10'h6) && 
                    |-------6--------|    |-------7--------|    |-------8--------|    |-------9--------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'h7) && (d[12:3] != 10'h8) && (d[12:3] != 10'h9) && (d[12:3] != 10'hA) && 
                    |-------10-------|    |-------11-------|    |-------12-------|    |-------13-------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hB) && (d[12:3] != 10'hC) && (d[12:3] != 10'hD) && (d[12:3] != 10'hE) && 
                    |-------14-------|    |-------15-------|    |-------16-------|    |-------17-------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hF) && (d[12:3] != 10'h10) && (d[12:3] != 10'h11) && (d[12:3] != 10'h12) && 
                    |-------18-------|    |-------19--------|    |-------20--------|    |-------21--------|    
                    ---------------------------------------------88---------------------------------------------
                    ---------------------------------------------89---------------------------------------------
                    --------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h13) && (d[12:3] != 10'h14) && (d[12:3] != 10'h15) && (d[12:3] != 10'h16) && 
                    |-------22--------|    |-------23--------|    |-------24--------|    |-------25--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h17) && (d[12:3] != 10'h18) && (d[12:3] != 10'h19) && (d[12:3] != 10'h1A) && 
                    |-------26--------|    |-------27--------|    |-------28--------|    |-------29--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1B) && (d[12:3] != 10'h1C) && (d[12:3] != 10'h1D) && (d[12:3] != 10'h1E) && 
                    |-------30--------|    |-------31--------|    |-------32--------|    |-------33--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1F) && (d[12:3] != 10'h20) && (d[12:3] != 10'h21) && (d[12:3] != 10'h22) && 
                    |-------34--------|    |-------35--------|    |-------36--------|    |-------37--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h23) && (d[12:3] != 10'h24) && (d[12:3] != 10'h25) && (d[12:3] != 10'h26) && 
                    |-------38--------|    |-------39--------|    |-------40--------|    |-------41--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h27) && (d[12:3] != 10'h28) && (d[12:3] != 10'h29) && (d[12:3] != 10'h2A) && 
                    |-------42--------|    |-------43--------|    |-------44--------|    |-------45--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2B) && (d[12:3] != 10'h2C) && (d[12:3] != 10'h2D) && (d[12:3] != 10'h2E) && 
                    |-------46--------|    |-------47--------|    |-------48--------|    |-------49--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2F) && (d[12:3] != 10'h30) && (d[12:3] != 10'h31) && (d[12:3] != 10'h32) && 
                    |-------50--------|    |-------51--------|    |-------52--------|    |-------53--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h33) && (d[12:3] != 10'h34) && (d[12:3] != 10'h35) && (d[12:3] != 10'h36) && 
                    |-------54--------|    |-------55--------|    |-------56--------|    |-------57--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h37) && (d[12:3] != 10'h38) && (d[12:3] != 10'h39) && (d[12:3] != 10'h3A) && 
                    |-------58--------|    |-------59--------|    |-------60--------|    |-------61--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3B) && (d[12:3] != 10'h3C) && (d[12:3] != 10'h3D) && (d[12:3] != 10'h3E) && 
                    |-------62--------|    |-------63--------|    |-------64--------|    |-------65--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3F) && (d[12:3] != 10'h40) && (d[12:3] != 10'h41) && (d[12:3] != 10'h42) && 
                    |-------66--------|    |-------67--------|    |-------68--------|    |-------69--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h43) && (d[12:3] != 10'h44) && (d[12:3] != 10'h45) && (d[12:3] != 10'h46) && 
                    |-------70--------|    |-------71--------|    |-------72--------|    |-------73--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h47) && (d[12:3] != 10'h48) && (d[12:3] != 10'h49) && (d[12:3] != 10'h4A) && 
                    |-------74--------|    |-------75--------|    |-------76--------|    |-------77--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4B) && (d[12:3] != 10'h4C) && (d[12:3] != 10'h4D) && (d[12:3] != 10'h4E) && 
                    |-------78--------|    |-------79--------|    |-------80--------|    |-------81--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4F) && (d[12:3] != 10'h50) && (d[12:3] != 10'h51) && (d[12:3] != 10'h52) && 
                    |-------82--------|    |-------83--------|    |-------84--------|    |-------85--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h53) && (d[12:3] != 10'h54))) | 
                    |-------86--------|    |-------87--------|     
                    --------------------88--------------------|    
                    ---------------------89--------------------|   
                    ----------------------169-----------------------
                    ( e  & ((d[27:16] == 12'h0) && (d[12:3] != 10'h0) && (d[12:3] != 10'h1) && (d[12:3] != 10'h2) && 
                            |-------90--------|    |-------91-------|    |-------92-------|    |-------93-------|    
                           |-------------------------------------------167--------------------------------------------
                    |----------------------------------------------168------------------------------------------------
                    -----------------------------------------------169------------------------------------------------
                    (d[12:3] != 10'h3) && (d[12:3] != 10'h4) && (d[12:3] != 10'h5) && (d[12:3] != 10'h6) && 
                    |-------94-------|    |-------95-------|    |-------96-------|    |-------97-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'h7) && (d[12:3] != 10'h8) && (d[12:3] != 10'h9) && (d[12:3] != 10'hA) && 
                    |-------98-------|    |-------99-------|    |------100-------|    |------101-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hB) && (d[12:3] != 10'hC) && (d[12:3] != 10'hD) && (d[12:3] != 10'hE) && 
                    |------102-------|    |------103-------|    |------104-------|    |------105-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hF) && (d[12:3] != 10'h10) && (d[12:3] != 10'h11) && (d[12:3] != 10'h12) && 
                    |------106-------|    |-------107-------|    |-------108-------|    |-------109-------|    
                    --------------------------------------------167---------------------------------------------
                    --------------------------------------------168---------------------------------------------
                    --------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h13) && (d[12:3] != 10'h14) && (d[12:3] != 10'h15) && (d[12:3] != 10'h16) && 
                    |-------110-------|    |-------111-------|    |-------112-------|    |-------113-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h17) && (d[12:3] != 10'h18) && (d[12:3] != 10'h19) && (d[12:3] != 10'h1A) && 
                    |-------114-------|    |-------115-------|    |-------116-------|    |-------117-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1B) && (d[12:3] != 10'h1C) && (d[12:3] != 10'h1D) && (d[12:3] != 10'h1E) && 
                    |-------118-------|    |-------119-------|    |-------120-------|    |-------121-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1F) && (d[12:3] != 10'h20) && (d[12:3] != 10'h21) && (d[12:3] != 10'h22) && 
                    |-------122-------|    |-------123-------|    |-------124-------|    |-------125-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h23) && (d[12:3] != 10'h24) && (d[12:3] != 10'h25) && (d[12:3] != 10'h26) && 
                    |-------126-------|    |-------127-------|    |-------128-------|    |-------129-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h27) && (d[12:3] != 10'h28) && (d[12:3] != 10'h29) && (d[12:3] != 10'h2A) && 
                    |-------130-------|    |-------131-------|    |-------132-------|    |-------133-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2B) && (d[12:3] != 10'h2C) && (d[12:3] != 10'h2D) && (d[12:3] != 10'h2E) && 
                    |-------134-------|    |-------135-------|    |-------136-------|    |-------137-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2F) && (d[12:3] != 10'h30) && (d[12:3] != 10'h31) && (d[12:3] != 10'h32) && 
                    |-------138-------|    |-------139-------|    |-------140-------|    |-------141-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h33) && (d[12:3] != 10'h34) && (d[12:3] != 10'h35) && (d[12:3] != 10'h36) && 
                    |-------142-------|    |-------143-------|    |-------144-------|    |-------145-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h37) && (d[12:3] != 10'h38) && (d[12:3] != 10'h39) && (d[12:3] != 10'h3A) && 
                    |-------146-------|    |-------147-------|    |-------148-------|    |-------149-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3B) && (d[12:3] != 10'h3C) && (d[12:3] != 10'h3D) && (d[12:3] != 10'h3E) && 
                    |-------150-------|    |-------151-------|    |-------152-------|    |-------153-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3F) && (d[12:3] != 10'h40) && (d[12:3] != 10'h41) && (d[12:3] != 10'h42) && 
                    |-------154-------|    |-------155-------|    |-------156-------|    |-------157-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h43) && (d[12:3] != 10'h44) && (d[12:3] != 10'h45) && (d[12:3] != 10'h46) && 
                    |-------158-------|    |-------159-------|    |-------160-------|    |-------161-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h47) && (d[12:3] != 10'h48) && (d[12:3] != 10'h49) && (d[12:3] != 10'h4A) && 
                    |-------162-------|    |-------163-------|    |-------164-------|    |-------165-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4B))))
                    |-------166-------|   
                    --------167--------|  
                    ---------168--------| 
                    ---------169---------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 3   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
             *

        Expression 4   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 5   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 6   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 7   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 8   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 9   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 10   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 11   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 12   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 13   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 14   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 15   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 16   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 17   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 18   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 19   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 20   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 21   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 22   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 23   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 24   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 25   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 26   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 27   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 28   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 29   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 30   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 31   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 32   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 33   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 34   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 35   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 36   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 37   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 38   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 39   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 40   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 41   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 42   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 43   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 44   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 45   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 46   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 47   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 48   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 49   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 50   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 51   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 52   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 53   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 54   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 55   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 56   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 57   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 58   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 59   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 60   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 61   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 62   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 63   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 64   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 65   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 66   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 67   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 68   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 69   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 70   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 71   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 72   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 73   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 74   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 75   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 76   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 77   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 78   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 79   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 80   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 81   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 82   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 83   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 84   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 85   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 86   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 87   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 88   (1/87)
        ^^^^^^^^^^^^^ - &&
         2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 | 16 | 17 | 18 | 19 | 20 | 21 | 22 | 23 | 24 |
        =0=|=0=|=0=|=0=|=0=|=0=|=0=|=0=|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *       *   *   *   *   *   *   *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         25 | 26 | 27 | 28 | 29 | 30 | 31 | 32 | 33 | 34 | 35 | 36 | 37 | 38 | 39 | 40 | 41 | 42 | 43 | 44 | 45 | 46 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         47 | 48 | 49 | 50 | 51 | 52 | 53 | 54 | 55 | 56 | 57 | 58 | 59 | 60 | 61 | 62 | 63 | 64 | 65 | 66 | 67 | 68 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         69 | 70 | 71 | 72 | 73 | 74 | 75 | 76 | 77 | 78 | 79 | 80 | 81 | 82 | 83 | 84 | 85 | 86 | 87 | All
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|==1==
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *     *  

        Expression 89   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 90   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 91   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
             *

        Expression 92   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 93   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 94   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 95   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 96   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 97   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 98   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 99   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 100   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 101   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 102   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 103   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 104   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 105   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 106   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 107   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 108   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 109   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 110   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 111   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 112   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 113   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 114   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 115   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 116   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 117   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 118   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 119   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 120   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 121   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 122   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 123   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 124   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 125   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 126   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 127   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 128   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 129   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 130   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 131   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 132   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 133   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 134   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 135   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 136   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 137   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 138   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 139   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 140   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 141   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 142   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 143   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 144   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 145   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 146   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 147   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 148   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 149   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 150   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 151   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 152   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 153   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 154   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 155   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 156   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 157   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 158   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 159   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 160   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 161   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 162   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 163   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 164   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 165   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 166   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 167   (1/78)
        ^^^^^^^^^^^^^ - &&
         90 | 91 | 92 | 93 | 94 | 95 | 96 | 97 | 98 | 99 | 100 | 101 | 102 | 103 | 104 | 105 | 106 | 107 | 108 | 109 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *         *    *    *    *    *    *    *    *    *     *     *     *     *     *     *     *     *     *    

         110 | 111 | 112 | 113 | 114 | 115 | 116 | 117 | 118 | 119 | 120 | 121 | 122 | 123 | 124 | 125 | 126 | 127 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         128 | 129 | 130 | 131 | 132 | 133 | 134 | 135 | 136 | 137 | 138 | 139 | 140 | 141 | 142 | 143 | 144 | 145 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         146 | 147 | 148 | 149 | 150 | 151 | 152 | 153 | 154 | 155 | 156 | 157 | 158 | 159 | 160 | 161 | 162 | 163 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         164 | 165 | 166 | All
        =0===|=0===|=0===|==1==
         *     *     *      *  

        Expression 168   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 169   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp1.v               0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT long_exp1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : long_exp1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/    0/    1      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/   29/   29        0%             0/   29/   29        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 25'h000_0000
      ......................... 1->0: 25'h000_0000 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                           169/ 338/ 507       33%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              8:    assign  a  = ((( b  |  c ) & 
                                   |----1----|   
                                  |------89-------
                                 |------169-------
                    ((d[27:16] == 12'h0) && 
                     |--------2--------|    
                    |----------88------------
                    -----------89------------
                    -----------169-----------
                    (d[12:3] != 10'h0) && 
                    |-------3--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h1) && 
                    |-------4--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h2) && 
                    |-------5--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h3) && 
                    |-------6--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h4) && 
                    |-------7--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h5) && 
                    |-------8--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h6) && 
                    |-------9--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h7) && 
                    |-------10-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h8) && 
                    |-------11-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h9) && 
                    |-------12-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hA) && 
                    |-------13-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hB) && 
                    |-------14-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hC) && 
                    |-------15-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hD) && 
                    |-------16-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hE) && 
                    |-------17-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hF) && 
                    |-------18-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h10) && 
                    |-------19--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h11) && 
                    |-------20--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h12) && 
                    |-------21--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h13) && 
                    |-------22--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h14) && 
                    |-------23--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h15) && 
                    |-------24--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h16) && 
                    |-------25--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h17) && 
                    |-------26--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h18) && 
                    |-------27--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h19) && 
                    |-------28--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1A) && 
                    |-------29--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1B) && 
                    |-------30--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1C) && 
                    |-------31--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1D) && 
                    |-------32--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1E) && 
                    |-------33--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1F) && 
                    |-------34--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h20) && 
                    |-------35--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h21) && 
                    |-------36--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h22) && 
                    |-------37--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h23) && 
                    |-------38--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h24) && 
                    |-------39--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h25) && 
                    |-------40--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h26) && 
                    |-------41--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h27) && 
                    |-------42--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h28) && 
                    |-------43--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h29) && 
                    |-------44--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2A) && 
                    |-------45--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2B) && 
                    |-------46--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2C) && 
                    |-------47--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2D) && 
                    |-------48--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2E) && 
                    |-------49--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2F) && 
                    |-------50--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h30) && 
                    |-------51--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h31) && 
                    |-------52--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h32) && 
                    |-------53--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h33) && 
                    |-------54--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h34) && 
                    |-------55--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h35) && 
                    |-------56--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h36) && 
                    |-------57--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h37) && 
                    |-------58--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h38) && 
                    |-------59--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h39) && 
                    |-------60--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3A) && 
                    |-------61--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3B) && 
                    |-------62--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3C) && 
                    |-------63--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3D) && 
                    |-------64--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3E) && 
                    |-------65--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3F) && 
                    |-------66--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h40) && 
                    |-------67--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h41) && 
                    |-------68--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h42) && 
                    |-------69--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h43) && 
                    |-------70--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h44) && 
                    |-------71--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h45) && 
                    |-------72--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h46) && 
                    |-------73--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h47) && 
                    |-------74--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h48) && 
                    |-------75--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h49) && 
                    |-------76--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4A) && 
                    |-------77--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4B) && 
                    |-------78--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4C) && 
                    |-------79--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4D) && 
                    |-------80--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4E) && 
                    |-------81--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4F) && 
                    |-------82--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h50) && 
                    |-------83--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h51) && 
                    |-------84--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h52) && 
                    |-------85--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h53) && 
                    |-------86--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h54))) | 
                    |-------87--------|     
                    ---------88--------|    
                    ---------89---------|   
                    -----------169-----------
                    ( e  & 
                    |-168---
                    --169---
                    ((d[27:16] == 12'h0) && 
                     |-------90--------|    
                    |----------167-----------
                    -----------168-----------
                    -----------169-----------
                    (d[12:3] != 10'h0) && 
                    |-------91-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h1) && 
                    |-------92-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h2) && 
                    |-------93-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h3) && 
                    |-------94-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h4) && 
                    |-------95-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h5) && 
                    |-------96-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h6) && 
                    |-------97-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h7) && 
                    |-------98-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h8) && 
                    |-------99-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h9) && 
                    |------100-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hA) && 
                    |------101-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hB) && 
                    |------102-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hC) && 
                    |------103-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hD) && 
                    |------104-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hE) && 
                    |------105-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hF) && 
                    |------106-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h10) && 
                    |-------107-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h11) && 
                    |-------108-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h12) && 
                    |-------109-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h13) && 
                    |-------110-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h14) && 
                    |-------111-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h15) && 
                    |-------112-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h16) && 
                    |-------113-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h17) && 
                    |-------114-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h18) && 
                    |-------115-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h19) && 
                    |-------116-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1A) && 
                    |-------117-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1B) && 
                    |-------118-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1C) && 
                    |-------119-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1D) && 
                    |-------120-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1E) && 
                    |-------121-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1F) && 
                    |-------122-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h20) && 
                    |-------123-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h21) && 
                    |-------124-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h22) && 
                    |-------125-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h23) && 
                    |-------126-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h24) && 
                    |-------127-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h25) && 
                    |-------128-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h26) && 
                    |-------129-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h27) && 
                    |-------130-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h28) && 
                    |-------131-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h29) && 
                    |-------132-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2A) && 
                    |-------133-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2B) && 
                    |-------134-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2C) && 
                    |-------135-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2D) && 
                    |-------136-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2E) && 
                    |-------137-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2F) && 
                    |-------138-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h30) && 
                    |-------139-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h31) && 
                    |-------140-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h32) && 
                    |-------141-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h33) && 
                    |-------142-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h34) && 
                    |-------143-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h35) && 
                    |-------144-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h36) && 
                    |-------145-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h37) && 
                    |-------146-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h38) && 
                    |-------147-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h39) && 
                    |-------148-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3A) && 
                    |-------149-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3B) && 
                    |-------150-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3C) && 
                    |-------151-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3D) && 
                    |-------152-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3E) && 
                    |-------153-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3F) && 
                    |-------154-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h40) && 
                    |-------155-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h41) && 
                    |-------156-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h42) && 
                    |-------157-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h43) && 
                    |-------158-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h44) && 
                    |-------159-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h45) && 
                    |-------160-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h46) && 
                    |-------161-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h47) && 
                    |-------162-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h48) && 
                    |-------163-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h49) && 
                    |-------164-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h4A) && 
                    |-------165-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h4B))))
                    |-------166-------|   
                    --------167--------|  
                    ---------168--------| 
                    ---------169---------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 3   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
             *

        Expression 4   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 5   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 6   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 7   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 8   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 9   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 10   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 11   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 12   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 13   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 14   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 15   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 16   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 17   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 18   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 19   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 20   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 21   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 22   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 23   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 24   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 25   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 26   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 27   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 28   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 29   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 30   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 31   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 32   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 33   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 34   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 35   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 36   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 37   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 38   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 39   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 40   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 41   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 42   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 43   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 44   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 45   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 46   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 47   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 48   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 49   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 50   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 51   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 52   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 53   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 54   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 55   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 56   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 57   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 58   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 59   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 60   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 61   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 62   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 63   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 64   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 65   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 66   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 67   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 68   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 69   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 70   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 71   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 72   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 73   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 74   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 75   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 76   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 77   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 78   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 79   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 80   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 81   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 82   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 83   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 84   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 85   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 86   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 87   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 88   (1/87)
        ^^^^^^^^^^^^^ - &&
         2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 | 16 | 17 | 18 | 19 | 20 | 21 | 22 | 23 | 24 |
        =0=|=0=|=0=|=0=|=0=|=0=|=0=|=0=|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *       *   *   *   *   *   *   *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         25 | 26 | 27 | 28 | 29 | 30 | 31 | 32 | 33 | 34 | 35 | 36 | 37 | 38 | 39 | 40 | 41 | 42 | 43 | 44 | 45 | 46 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         47 | 48 | 49 | 50 | 51 | 52 | 53 | 54 | 55 | 56 | 57 | 58 | 59 | 60 | 61 | 62 | 63 | 64 | 65 | 66 | 67 | 68 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         69 | 70 | 71 | 72 | 73 | 74 | 75 | 76 | 77 | 78 | 79 | 80 | 81 | 82 | 83 | 84 | 85 | 86 | 87 | All
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|==1==
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *     *  

        Expression 89   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 90   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 91   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
             *

        Expression 92   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 93   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 94   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 95   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 96   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 97   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 98   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 99   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 100   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 101   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 102   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 103   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 104   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 105   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 106   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 107   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 108   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 109   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 110   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 111   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 112   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 113   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 114   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 115   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 116   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 117   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 118   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 119   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 120   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 121   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 122   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 123   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 124   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 125   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 126   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 127   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 128   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 129   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 130   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 131   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 132   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 133   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 134   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 135   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 136   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 137   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 138   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 139   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 140   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 141   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 142   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 143   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 144   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 145   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 146   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 147   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 148   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 149   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 150   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 151   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 152   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 153   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 154   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 155   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 156   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 157   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 158   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 159   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 160   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 161   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 162   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 163   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 164   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 165   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 166   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 167   (1/78)
        ^^^^^^^^^^^^^ - &&
         90 | 91 | 92 | 93 | 94 | 95 | 96 | 97 | 98 | 99 | 100 | 101 | 102 | 103 | 104 | 105 | 106 | 107 | 108 | 109 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *         *    *    *    *    *    *    *    *    *     *     *     *     *     *     *     *     *     *    

         110 | 111 | 112 | 113 | 114 | 115 | 116 | 117 | 118 | 119 | 120 | 121 | 122 | 123 | 124 | 125 | 126 | 127 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         128 | 129 | 130 | 131 | 132 | 133 | 134 | 135 | 136 | 137 | 138 | 139 | 140 | 141 | 142 | 143 | 144 | 145 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         146 | 147 | 148 | 149 | 150 | 151 | 152 | 153 | 154 | 155 | 156 | 157 | 158 | 159 | 160 | 161 | 162 | 163 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         164 | 165 | 166 | All
        =0===|=0===|=0===|==1==
         *     *     *      *  

        Expression 168   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 169   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT long_exp1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : long_exp1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/    0/    1      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/   29/   29        0%             0/   29/   29        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 25'h000_0000
      ......................... 1->0: 25'h000_0000 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                           169/ 338/ 507       33%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              8:    assign  a  = ((( b  |  c ) & 
                                   |----1----|   
                                  |------89-------
                                 |------169-------
                    ((d[27:16] == 12'h0) && (d[12:3] != 10'h0) && (d[12:3] != 10'h1) && (d[12:3] != 10'h2) && 
                     |--------2--------|    |-------3--------|    |-------4--------|    |-------5--------|    
                    |-------------------------------------------88---------------------------------------------
                    --------------------------------------------89---------------------------------------------
                    --------------------------------------------169--------------------------------------------
                    (d[12:3] != 10'h3) && (d[12:3] != 10'h4) && (d[12:3] != 10'h5) && (d[12:3] != 10'h6) && 
                    |-------6--------|    |-------7--------|    |-------8--------|    |-------9--------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'h7) && (d[12:3] != 10'h8) && (d[12:3] != 10'h9) && (d[12:3] != 10'hA) && 
                    |-------10-------|    |-------11-------|    |-------12-------|    |-------13-------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hB) && (d[12:3] != 10'hC) && (d[12:3] != 10'hD) && (d[12:3] != 10'hE) && 
                    |-------14-------|    |-------15-------|    |-------16-------|    |-------17-------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hF) && (d[12:3] != 10'h10) && (d[12:3] != 10'h11) && (d[12:3] != 10'h12) && 
                    |-------18-------|    |-------19--------|    |-------20--------|    |-------21--------|    
                    ---------------------------------------------88---------------------------------------------
                    ---------------------------------------------89---------------------------------------------
                    --------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h13) && (d[12:3] != 10'h14) && (d[12:3] != 10'h15) && (d[12:3] != 10'h16) && 
                    |-------22--------|    |-------23--------|    |-------24--------|    |-------25--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h17) && (d[12:3] != 10'h18) && (d[12:3] != 10'h19) && (d[12:3] != 10'h1A) && 
                    |-------26--------|    |-------27--------|    |-------28--------|    |-------29--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1B) && (d[12:3] != 10'h1C) && (d[12:3] != 10'h1D) && (d[12:3] != 10'h1E) && 
                    |-------30--------|    |-------31--------|    |-------32--------|    |-------33--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1F) && (d[12:3] != 10'h20) && (d[12:3] != 10'h21) && (d[12:3] != 10'h22) && 
                    |-------34--------|    |-------35--------|    |-------36--------|    |-------37--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h23) && (d[12:3] != 10'h24) && (d[12:3] != 10'h25) && (d[12:3] != 10'h26) && 
                    |-------38--------|    |-------39--------|    |-------40--------|    |-------41--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h27) && (d[12:3] != 10'h28) && (d[12:3] != 10'h29) && (d[12:3] != 10'h2A) && 
                    |-------42--------|    |-------43--------|    |-------44--------|    |-------45--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2B) && (d[12:3] != 10'h2C) && (d[12:3] != 10'h2D) && (d[12:3] != 10'h2E) && 
                    |-------46--------|    |-------47--------|    |-------48--------|    |-------49--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2F) && (d[12:3] != 10'h30) && (d[12:3] != 10'h31) && (d[12:3] != 10'h32) && 
                    |-------50--------|    |-------51--------|    |-------52--------|    |-------53--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h33) && (d[12:3] != 10'h34) && (d[12:3] != 10'h35) && (d[12:3] != 10'h36) && 
                    |-------54--------|    |-------55--------|    |-------56--------|    |-------57--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h37) && (d[12:3] != 10'h38) && (d[12:3] != 10'h39) && (d[12:3] != 10'h3A) && 
                    |-------58--------|    |-------59--------|    |-------60--------|    |-------61--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3B) && (d[12:3] != 10'h3C) && (d[12:3] != 10'h3D) && (d[12:3] != 10'h3E) && 
                    |-------62--------|    |-------63--------|    |-------64--------|    |-------65--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3F) && (d[12:3] != 10'h40) && (d[12:3] != 10'h41) && (d[12:3] != 10'h42) && 
                    |-------66--------|    |-------67--------|    |-------68--------|    |-------69--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h43) && (d[12:3] != 10'h44) && (d[12:3] != 10'h45) && (d[12:3] != 10'h46) && 
                    |-------70--------|    |-------71--------|    |-------72--------|    |-------73--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h47) && (d[12:3] != 10'h48) && (d[12:3] != 10'h49) && (d[12:3] != 10'h4A) && 
                    |-------74--------|    |-------75--------|    |-------76--------|    |-------77--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4B) && (d[12:3] != 10'h4C) && (d[12:3] != 10'h4D) && (d[12:3] != 10'h4E) && 
                    |-------78--------|    |-------79--------|    |-------80--------|    |-------81--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4F) && (d[12:3] != 10'h50) && (d[12:3] != 10'h51) && (d[12:3] != 10'h52) && 
                    |-------82--------|    |-------83--------|    |-------84--------|    |-------85--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h53) && (d[12:3] != 10'h54))) | 
                    |-------86--------|    |-------87--------|     
                    --------------------88--------------------|    
                    ---------------------89--------------------|   
                    ----------------------169-----------------------
                    ( e  & ((d[27:16] == 12'h0) && (d[12:3] != 10'h0) && (d[12:3] != 10'h1) && (d[12:3] != 10'h2) && 
                            |-------90--------|    |-------91-------|    |-------92-------|    |-------93-------|    
                           |-------------------------------------------167--------------------------------------------
                    |----------------------------------------------168------------------------------------------------
                    -----------------------------------------------169------------------------------------------------
                    (d[12:3] != 10'h3) && (d[12:3] != 10'h4) && (d[12:3] != 10'h5) && (d[12:3] != 10'h6) && 
                    |-------94-------|    |-------95-------|    |-------96-------|    |-------97-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'h7) && (d[12:3] != 10'h8) && (d[12:3] != 10'h9) && (d[12:3] != 10'hA) && 
                    |-------98-------|    |-------99-------|    |------100-------|    |------101-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hB) && (d[12:3] != 10'hC) && (d[12:3] != 10'hD) && (d[12:3] != 10'hE) && 
                    |------102-------|    |------103-------|    |------104-------|    |------105-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hF) && (d[12:3] != 10'h10) && (d[12:3] != 10'h11) && (d[12:3] != 10'h12) && 
                    |------106-------|    |-------107-------|    |-------108-------|    |-------109-------|    
                    --------------------------------------------167---------------------------------------------
                    --------------------------------------------168---------------------------------------------
                    --------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h13) && (d[12:3] != 10'h14) && (d[12:3] != 10'h15) && (d[12:3] != 10'h16) && 
                    |-------110-------|    |-------111-------|    |-------112-------|    |-------113-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h17) && (d[12:3] != 10'h18) && (d[12:3] != 10'h19) && (d[12:3] != 10'h1A) && 
                    |-------114-------|    |-------115-------|    |-------116-------|    |-------117-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1B) && (d[12:3] != 10'h1C) && (d[12:3] != 10'h1D) && (d[12:3] != 10'h1E) && 
                    |-------118-------|    |-------119-------|    |-------120-------|    |-------121-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1F) && (d[12:3] != 10'h20) && (d[12:3] != 10'h21) && (d[12:3] != 10'h22) && 
                    |-------122-------|    |-------123-------|    |-------124-------|    |-------125-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h23) && (d[12:3] != 10'h24) && (d[12:3] != 10'h25) && (d[12:3] != 10'h26) && 
                    |-------126-------|    |-------127-------|    |-------128-------|    |-------129-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h27) && (d[12:3] != 10'h28) && (d[12:3] != 10'h29) && (d[12:3] != 10'h2A) && 
                    |-------130-------|    |-------131-------|    |-------132-------|    |-------133-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2B) && (d[12:3] != 10'h2C) && (d[12:3] != 10'h2D) && (d[12:3] != 10'h2E) && 
                    |-------134-------|    |-------135-------|    |-------136-------|    |-------137-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2F) && (d[12:3] != 10'h30) && (d[12:3] != 10'h31) && (d[12:3] != 10'h32) && 
                    |-------138-------|    |-------139-------|    |-------140-------|    |-------141-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h33) && (d[12:3] != 10'h34) && (d[12:3] != 10'h35) && (d[12:3] != 10'h36) && 
                    |-------142-------|    |-------143-------|    |-------144-------|    |-------145-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h37) && (d[12:3] != 10'h38) && (d[12:3] != 10'h39) && (d[12:3] != 10'h3A) && 
                    |-------146-------|    |-------147-------|    |-------148-------|    |-------149-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3B) && (d[12:3] != 10'h3C) && (d[12:3] != 10'h3D) && (d[12:3] != 10'h3E) && 
                    |-------150-------|    |-------151-------|    |-------152-------|    |-------153-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3F) && (d[12:3] != 10'h40) && (d[12:3] != 10'h41) && (d[12:3] != 10'h42) && 
                    |-------154-------|    |-------155-------|    |-------156-------|    |-------157-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h43) && (d[12:3] != 10'h44) && (d[12:3] != 10'h45) && (d[12:3] != 10'h46) && 
                    |-------158-------|    |-------159-------|    |-------160-------|    |-------161-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h47) && (d[12:3] != 10'h48) && (d[12:3] != 10'h49) && (d[12:3] != 10'h4A) && 
                    |-------162-------|    |-------163-------|    |-------164-------|    |-------165-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4B))))
                    |-------166-------|   
                    --------167--------|  
                    ---------168--------| 
                    ---------169---------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 3   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
             *

        Expression 4   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 5   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 6   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 7   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 8   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 9   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 10   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 11   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 12   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 13   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 14   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 15   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 16   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 17   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 18   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 19   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 20   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 21   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 22   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 23   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 24   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 25   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 26   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 27   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 28   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 29   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 30   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 31   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 32   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 33   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 34   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 35   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 36   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 37   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 38   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 39   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 40   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 41   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 42   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 43   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 44   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 45   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 46   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 47   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 48   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 49   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 50   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 51   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 52   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 53   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 54   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 55   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 56   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 57   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 58   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 59   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 60   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 61   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 62   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 63   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 64   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 65   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 66   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 67   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 68   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 69   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 70   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 71   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 72   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 73   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 74   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 75   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 76   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 77   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 78   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 79   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 80   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 81   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 82   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 83   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 84   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 85   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 86   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 87   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 88   (1/87)
        ^^^^^^^^^^^^^ - &&
         2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 | 16 | 17 | 18 | 19 | 20 | 21 | 22 | 23 | 24 |
        =0=|=0=|=0=|=0=|=0=|=0=|=0=|=0=|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *       *   *   *   *   *   *   *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         25 | 26 | 27 | 28 | 29 | 30 | 31 | 32 | 33 | 34 | 35 | 36 | 37 | 38 | 39 | 40 | 41 | 42 | 43 | 44 | 45 | 46 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         47 | 48 | 49 | 50 | 51 | 52 | 53 | 54 | 55 | 56 | 57 | 58 | 59 | 60 | 61 | 62 | 63 | 64 | 65 | 66 | 67 | 68 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         69 | 70 | 71 | 72 | 73 | 74 | 75 | 76 | 77 | 78 | 79 | 80 | 81 | 82 | 83 | 84 | 85 | 86 | 87 | All
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|==1==
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *     *  

        Expression 89   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 90   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 91   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
             *

        Expression 92   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 93   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 94   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 95   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 96   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 97   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 98   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 99   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 100   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 101   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 102   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 103   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 104   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 105   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 106   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 107   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 108   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 109   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 110   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 111   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 112   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 113   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 114   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 115   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 116   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 117   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 118   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 119   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 120   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 121   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 122   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 123   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 124   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 125   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 126   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 127   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 128   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 129   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 130   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 131   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 132   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 133   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 134   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 135   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 136   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 137   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 138   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 139   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 140   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 141   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 142   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 143   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 144   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 145   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 146   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 147   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 148   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 149   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 150   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 151   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 152   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 153   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 154   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 155   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 156   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 157   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 158   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 159   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 160   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 161   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 162   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 163   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 164   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 165   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 166   (1/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *    

        Expression 167   (1/78)
        ^^^^^^^^^^^^^ - &&
         90 | 91 | 92 | 93 | 94 | 95 | 96 | 97 | 98 | 99 | 100 | 101 | 102 | 103 | 104 | 105 | 106 | 107 | 108 | 109 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *         *    *    *    *    *    *    *    *    *     *     *     *     *     *     *     *     *     *    

         110 | 111 | 112 | 113 | 114 | 115 | 116 | 117 | 118 | 119 | 120 | 121 | 122 | 123 | 124 | 125 | 126 | 127 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         128 | 129 | 130 | 131 | 132 | 133 | 134 | 135 | 136 | 137 | 138 | 139 | 140 | 141 | 142 | 143 | 144 | 145 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         146 | 147 | 148 | 149 | 150 | 151 | 152 | 153 | 154 | 155 | 156 | 157 | 158 | 159 | 160 | 161 | 162 | 163 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         164 | 165 | 166 | All
        =0===|=0===|=0===|==1==
         *     *     *      *  

        Expression 168   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 169   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
