module main;

foo f();

endmodule

//-------------------------

module foo (
  a
);

output reg a;

endmodule
