module main;

foo #(2)       a();
foo #(3,4)     b();
foo #(.car(6)) c();

initial begin
        $dumpfile( "param10.5.vcd" );
        $dumpvars( 0, main );
        #10;
        $finish;
end

endmodule


module foo;

parameter bar = 1;

wire [(bar-1):0] b;
reg  [31:0]      c;

initial begin : foo_begin
	parameter car = 5;
	reg [(car-1):0] a;
	a = 1'b0;
end

initial begin
        c = 0;
        c = bar;
end

endmodule

/* HEADER
GROUPS param10.5 all iv vcs vcd lxt
SIM    param10.5 all iv vcd  : iverilog param10.5.v; ./a.out                             : param10.5.vcd
SIM    param10.5 all iv lxt  : iverilog param10.5.v; ./a.out -lxt2; mv param10.5.vcd param10.5.lxt : param10.5.lxt
SIM    param10.5 all vcs vcd : vcs +v2k param10.5.v; ./simv                                        : param10.5.vcd
SCORE  param10.5.vcd     : -t main -vcd param10.5.vcd -o param10.5.cdd -v param10.5.v : param10.5.cdd
SCORE  param10.5.lxt     : -t main -lxt param10.5.lxt -o param10.5.cdd -v param10.5.v : param10.5.cdd
REPORT param10.5.cdd 1   : -d v -o param10.5.rptM param10.5.cdd                         : param10.5.rptM
REPORT param10.5.cdd 2   : -d v -w -o param10.5.rptWM param10.5.cdd                     : param10.5.rptWM
REPORT param10.5.cdd 3   : -d v -i -o param10.5.rptI param10.5.cdd                      : param10.5.rptI
REPORT param10.5.cdd 4   : -d v -w -i -o param10.5.rptWI param10.5.cdd                  : param10.5.rptWI
*/

/* OUTPUT param10.5.cdd
5 1 * 6 0 0 0 0
3 0 main main param10.5.v 1 14
1 #car 0 0 0 32 0 14 0 0 0 0 0 0 0
3 0 foo main.a param10.5.v 17 35
2 1 24 8000c 2 3d 2100a 0 0 1 0 2 foo_begin
2 2 31 c000c 1 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 3 31 80008 0 1 400 0 0 c
2 4 31 8000c 1 37 1006 2 3
2 5 32 c000e 1 32 8 0 0 #bar
2 6 32 80008 0 1 400 0 0 c
2 7 32 8000e 1 37 a 5 6
1 #bar 0 0 0 32 0 4 0 0 0 0 0 0 0
1 b 0 21 30011 2 0 a
1 c 0 22 30011 32 16 2aa aa aa aa aa aa aa aa
4 1 0 0
4 7 0 0
4 4 7 7
3 1 foo.foo_begin main.a.foo_begin param10.5.v 24 28
2 8 27 50008 1 0 20004 0 0 1 1 0
2 9 27 10001 0 1 400 0 0 a
2 10 27 10008 1 37 11006 8 9
1 #car 0 0 0 32 0 11 0 0 0 0 0 0 0
1 a 0 26 30011 5 16 aa 2
4 10 0 0
3 0 foo main.b param10.5.v 17 35
2 11 24 8000c 2 3d 2100a 0 0 1 0 2 foo_begin
2 12 31 c000c 1 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 13 31 80008 0 1 400 0 0 c
2 14 31 8000c 1 37 1006 12 13
2 15 32 c000e 1 32 8 0 0 #bar
2 16 32 80008 0 1 400 0 0 c
2 17 32 8000e 1 37 a 15 16
1 #bar 0 0 0 32 0 5 0 0 0 0 0 0 0
1 b 0 21 30011 3 0 2a
1 c 0 22 30011 32 16 3aa aa aa aa aa aa aa aa
4 11 0 0
4 17 0 0
4 14 17 17
3 1 foo.foo_begin main.b.foo_begin param10.5.v 24 28
2 18 27 50008 1 0 20004 0 0 1 1 0
2 19 27 10001 0 1 400 0 0 a
2 20 27 10008 1 37 11006 18 19
1 #car 0 0 0 32 0 10 0 0 0 0 0 0 0
1 a 0 26 30011 4 16 aa
4 20 0 0
3 0 foo main.c param10.5.v 17 35
2 21 24 8000c 2 3d 2100a 0 0 1 0 2 foo_begin
2 22 31 c000c 1 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 23 31 80008 0 1 400 0 0 c
2 24 31 8000c 1 37 1006 22 23
2 25 32 c000e 1 32 8 0 0 #bar
2 26 32 80008 0 1 400 0 0 c
2 27 32 8000e 1 37 a 25 26
1 #bar 0 0 0 32 0 1 0 0 0 0 0 0 0
1 b 0 21 30011 1 0 2
1 c 0 22 30011 32 16 1aa aa aa aa aa aa aa aa
4 21 0 0
4 27 0 0
4 24 27 27
3 1 foo.foo_begin main.c.foo_begin param10.5.v 24 28
2 28 27 50008 1 0 20004 0 0 1 1 0
2 29 27 10001 0 1 400 0 0 a
2 30 27 10008 1 37 11006 28 29
1 #car 0 0 0 32 0 14 0 0 0 0 0 0 0
1 a 0 26 30011 6 16 aa a
4 30 0 0
*/

/* OUTPUT param10.5.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : param10.5.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    param10.5.v                0/    0/    0      100%
  foo                     param10.5.v                2/    0/    2      100%
  foo.foo_begin           param10.5.v                1/    0/    1      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    param10.5.v                0/    0/    0      100%             0/    0/    0      100%
  foo                     param10.5.v                2/   32/   34        6%             0/   34/   34        0%
  foo.foo_begin           param10.5.v                0/    5/    5        0%             0/    5/    5        0%
---------------------------------------------------------------------------------------------------------------------

    Module: foo, File: param10.5.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      b                         0->1: 2'h0
      ......................... 1->0: 2'h0 ...
      c                         0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0000 ...

    Named Block: foo.foo_begin, File: param10.5.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 5'h00
      ......................... 1->0: 5'h00 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              param10.5.v                         0/   0/   0      100%
  foo                               param10.5.v                         0/   0/   0      100%
  foo.foo_begin                     param10.5.v                         0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    param10.5.v               0/   0/   0      100%            0/   0/   0      100%
  foo                     param10.5.v               0/   0/   0      100%            0/   0/   0      100%
  foo.foo_begin           param10.5.v               0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT param10.5.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : param10.5.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    param10.5.v                0/    0/    0      100%
  foo                     param10.5.v                2/    0/    2      100%
  foo.foo_begin           param10.5.v                1/    0/    1      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    param10.5.v                0/    0/    0      100%             0/    0/    0      100%
  foo                     param10.5.v                2/   32/   34        6%             0/   34/   34        0%
  foo.foo_begin           param10.5.v                0/    5/    5        0%             0/    5/    5        0%
---------------------------------------------------------------------------------------------------------------------

    Module: foo, File: param10.5.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      b                         0->1: 2'h0
      ......................... 1->0: 2'h0 ...
      c                         0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0000 ...

    Named Block: foo.foo_begin, File: param10.5.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 5'h00
      ......................... 1->0: 5'h00 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              param10.5.v                         0/   0/   0      100%
  foo                               param10.5.v                         0/   0/   0      100%
  foo.foo_begin                     param10.5.v                         0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    param10.5.v               0/   0/   0      100%            0/   0/   0      100%
  foo                     param10.5.v               0/   0/   0      100%            0/   0/   0      100%
  foo.foo_begin           param10.5.v               0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT param10.5.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : param10.5.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%
  <NA>.main.a                                        2/    0/    2      100%
  <NA>.main.a.foo_begin                              1/    0/    1      100%
  <NA>.main.b                                        2/    0/    2      100%
  <NA>.main.b.foo_begin                              1/    0/    1      100%
  <NA>.main.c                                        2/    0/    2      100%
  <NA>.main.c.foo_begin                              1/    0/    1      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%             0/    0/    0      100%
  <NA>.main.a                                        1/   33/   34        3%             0/   34/   34        0%
  <NA>.main.a.foo_begin                              0/    5/    5        0%             0/    5/    5        0%
  <NA>.main.b                                        2/   33/   35        6%             0/   35/   35        0%
  <NA>.main.b.foo_begin                              0/    4/    4        0%             0/    4/    4        0%
  <NA>.main.c                                        1/   32/   33        3%             0/   33/   33        0%
  <NA>.main.c.foo_begin                              0/    6/    6        0%             0/    6/    6        0%
---------------------------------------------------------------------------------------------------------------------

    Module: foo, File: param10.5.v, Instance: <NA>.main.a
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      b                         0->1: 2'h0
      ......................... 1->0: 2'h0 ...
      c                         0->1: 32'h0000_0002
      ......................... 1->0: 32'h0000_0000 ...

    Named Block: foo.foo_begin, File: param10.5.v, Instance: <NA>.main.a.foo_begin
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 5'h00
      ......................... 1->0: 5'h00 ...

    Module: foo, File: param10.5.v, Instance: <NA>.main.b
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      b                         0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      c                         0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0000 ...

    Named Block: foo.foo_begin, File: param10.5.v, Instance: <NA>.main.b.foo_begin
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h0
      ......................... 1->0: 4'h0 ...

    Module: foo, File: param10.5.v, Instance: <NA>.main.c
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0000 ...

    Named Block: foo.foo_begin, File: param10.5.v, Instance: <NA>.main.c.foo_begin
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 6'h00
      ......................... 1->0: 6'h00 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%
  <NA>.main.a                                                           0/   0/   0      100%
  <NA>.main.a.foo_begin                                                 0/   0/   0      100%
  <NA>.main.b                                                           0/   0/   0      100%
  <NA>.main.b.foo_begin                                                 0/   0/   0      100%
  <NA>.main.c                                                           0/   0/   0      100%
  <NA>.main.c.foo_begin                                                 0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.a                                       0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.a.foo_begin                             0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.b                                       0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.b.foo_begin                             0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.c                                       0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.c.foo_begin                             0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT param10.5.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : param10.5.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%
  <NA>.main.a                                        2/    0/    2      100%
  <NA>.main.a.foo_begin                              1/    0/    1      100%
  <NA>.main.b                                        2/    0/    2      100%
  <NA>.main.b.foo_begin                              1/    0/    1      100%
  <NA>.main.c                                        2/    0/    2      100%
  <NA>.main.c.foo_begin                              1/    0/    1      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%             0/    0/    0      100%
  <NA>.main.a                                        1/   33/   34        3%             0/   34/   34        0%
  <NA>.main.a.foo_begin                              0/    5/    5        0%             0/    5/    5        0%
  <NA>.main.b                                        2/   33/   35        6%             0/   35/   35        0%
  <NA>.main.b.foo_begin                              0/    4/    4        0%             0/    4/    4        0%
  <NA>.main.c                                        1/   32/   33        3%             0/   33/   33        0%
  <NA>.main.c.foo_begin                              0/    6/    6        0%             0/    6/    6        0%
---------------------------------------------------------------------------------------------------------------------

    Module: foo, File: param10.5.v, Instance: <NA>.main.a
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      b                         0->1: 2'h0
      ......................... 1->0: 2'h0 ...
      c                         0->1: 32'h0000_0002
      ......................... 1->0: 32'h0000_0000 ...

    Named Block: foo.foo_begin, File: param10.5.v, Instance: <NA>.main.a.foo_begin
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 5'h00
      ......................... 1->0: 5'h00 ...

    Module: foo, File: param10.5.v, Instance: <NA>.main.b
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      b                         0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      c                         0->1: 32'h0000_0003
      ......................... 1->0: 32'h0000_0000 ...

    Named Block: foo.foo_begin, File: param10.5.v, Instance: <NA>.main.b.foo_begin
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h0
      ......................... 1->0: 4'h0 ...

    Module: foo, File: param10.5.v, Instance: <NA>.main.c
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 32'h0000_0001
      ......................... 1->0: 32'h0000_0000 ...

    Named Block: foo.foo_begin, File: param10.5.v, Instance: <NA>.main.c.foo_begin
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 6'h00
      ......................... 1->0: 6'h00 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%
  <NA>.main.a                                                           0/   0/   0      100%
  <NA>.main.a.foo_begin                                                 0/   0/   0      100%
  <NA>.main.b                                                           0/   0/   0      100%
  <NA>.main.b.foo_begin                                                 0/   0/   0      100%
  <NA>.main.c                                                           0/   0/   0      100%
  <NA>.main.c.foo_begin                                                 0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.a                                       0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.a.foo_begin                             0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.b                                       0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.b.foo_begin                             0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.c                                       0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.c.foo_begin                             0/   0/   0      100%            0/   0/   0      100%


*/
