module main;

reg         go;
reg         a;
reg         b, c;
reg  [27:3] d;
reg         e;

always @(posedge go)
  begin
   a <= (b | c) &
         ((d[27:16]==12'h0) &&
         (d[12:3] != 10'h000) &&
         (d[12:3] != 10'h001) &&
         (d[12:3] != 10'h002) &&
         (d[12:3] != 10'h003) &&
         (d[12:3] != 10'h004) &&
         (d[12:3] != 10'h005) &&
         (d[12:3] != 10'h006) &&
         (d[12:3] != 10'h007) &&
         (d[12:3] != 10'h008) &&
         (d[12:3] != 10'h009) &&
         (d[12:3] != 10'h00A) &&
         (d[12:3] != 10'h00B) &&
         (d[12:3] != 10'h00C) &&
         (d[12:3] != 10'h00D) &&
         (d[12:3] != 10'h00E) &&
         (d[12:3] != 10'h00F) &&
         (d[12:3] != 10'h010) &&
         (d[12:3] != 10'h011) &&
         (d[12:3] != 10'h012) &&
         (d[12:3] != 10'h013) &&
         (d[12:3] != 10'h014) &&
         (d[12:3] != 10'h015) &&
         (d[12:3] != 10'h016) &&
         (d[12:3] != 10'h017) &&
         (d[12:3] != 10'h018) &&
         (d[12:3] != 10'h019) &&
         (d[12:3] != 10'h01A) &&
         (d[12:3] != 10'h01B) &&
         (d[12:3] != 10'h01C) &&
         (d[12:3] != 10'h01D) &&
         (d[12:3] != 10'h01E) &&
         (d[12:3] != 10'h01F) &&
         (d[12:3] != 10'h020) &&
         (d[12:3] != 10'h021) &&
         (d[12:3] != 10'h022) &&
         (d[12:3] != 10'h023) &&
         (d[12:3] != 10'h024) &&
         (d[12:3] != 10'h025) &&
         (d[12:3] != 10'h026) &&
         (d[12:3] != 10'h027) &&
         (d[12:3] != 10'h028) &&
         (d[12:3] != 10'h029) &&
         (d[12:3] != 10'h02A) &&
         (d[12:3] != 10'h02B) &&
         (d[12:3] != 10'h02C) &&
         (d[12:3] != 10'h02D) &&
         (d[12:3] != 10'h02E) &&
         (d[12:3] != 10'h02F) &&
         (d[12:3] != 10'h030) &&
         (d[12:3] != 10'h031) &&
         (d[12:3] != 10'h032) &&
         (d[12:3] != 10'h033) &&
         (d[12:3] != 10'h034) &&
         (d[12:3] != 10'h035) &&
         (d[12:3] != 10'h036) &&
         (d[12:3] != 10'h037) &&
         (d[12:3] != 10'h038) &&
         (d[12:3] != 10'h039) &&
         (d[12:3] != 10'h03A) &&
         (d[12:3] != 10'h03B) &&
         (d[12:3] != 10'h03C) &&
         (d[12:3] != 10'h03D) &&
         (d[12:3] != 10'h03E) &&
         (d[12:3] != 10'h03F) &&
         (d[12:3] != 10'h040) &&
         (d[12:3] != 10'h041) &&
         (d[12:3] != 10'h042) &&
         (d[12:3] != 10'h043) &&
         (d[12:3] != 10'h044) &&
         (d[12:3] != 10'h045) &&
         (d[12:3] != 10'h046) &&
         (d[12:3] != 10'h047) &&
         (d[12:3] != 10'h048) &&
         (d[12:3] != 10'h049) &&
         (d[12:3] != 10'h04A) &&
         (d[12:3] != 10'h04B) &&
         (d[12:3] != 10'h04C) &&
         (d[12:3] != 10'h04D) &&
         (d[12:3] != 10'h04E) &&
         (d[12:3] != 10'h04F) &&
         (d[12:3] != 10'h050) &&
         (d[12:3] != 10'h051) &&
         (d[12:3] != 10'h052) &&
         (d[12:3] != 10'h053) &&
         (d[12:3] != 10'h054)) |
        e &
        ((d[27:16]==12'h0) &&
         (d[12:3] != 10'h000) &&
         (d[12:3] != 10'h001) &&
         (d[12:3] != 10'h002) &&
         (d[12:3] != 10'h003) &&
         (d[12:3] != 10'h004) &&
         (d[12:3] != 10'h005) &&
         (d[12:3] != 10'h006) &&
         (d[12:3] != 10'h007) &&
         (d[12:3] != 10'h008) &&
         (d[12:3] != 10'h009) &&
         (d[12:3] != 10'h00A) &&
         (d[12:3] != 10'h00B) &&
         (d[12:3] != 10'h00C) &&
         (d[12:3] != 10'h00D) &&
         (d[12:3] != 10'h00E) &&
         (d[12:3] != 10'h00F) &&
         (d[12:3] != 10'h010) &&
         (d[12:3] != 10'h011) &&
         (d[12:3] != 10'h012) &&
         (d[12:3] != 10'h013) &&
         (d[12:3] != 10'h014) &&
         (d[12:3] != 10'h015) &&
         (d[12:3] != 10'h016) &&
         (d[12:3] != 10'h017) &&
         (d[12:3] != 10'h018) &&
         (d[12:3] != 10'h019) &&
         (d[12:3] != 10'h01A) &&
         (d[12:3] != 10'h01B) &&
         (d[12:3] != 10'h01C) &&
         (d[12:3] != 10'h01D) &&
         (d[12:3] != 10'h01E) &&
         (d[12:3] != 10'h01F) &&
         (d[12:3] != 10'h020) &&
         (d[12:3] != 10'h021) &&
         (d[12:3] != 10'h022) &&
         (d[12:3] != 10'h023) &&
         (d[12:3] != 10'h024) &&
         (d[12:3] != 10'h025) &&
         (d[12:3] != 10'h026) &&
         (d[12:3] != 10'h027) &&
         (d[12:3] != 10'h028) &&
         (d[12:3] != 10'h029) &&
         (d[12:3] != 10'h02A) &&
         (d[12:3] != 10'h02B) &&
         (d[12:3] != 10'h02C) &&
         (d[12:3] != 10'h02D) &&
         (d[12:3] != 10'h02E) &&
         (d[12:3] != 10'h02F) &&
         (d[12:3] != 10'h030) &&
         (d[12:3] != 10'h031) &&
         (d[12:3] != 10'h032) &&
         (d[12:3] != 10'h033) &&
         (d[12:3] != 10'h034) &&
         (d[12:3] != 10'h035) &&
         (d[12:3] != 10'h036) &&
         (d[12:3] != 10'h037) &&
         (d[12:3] != 10'h038) &&
         (d[12:3] != 10'h039) &&
         (d[12:3] != 10'h03A) &&
         (d[12:3] != 10'h03B) &&
         (d[12:3] != 10'h03C) &&
         (d[12:3] != 10'h03D) &&
         (d[12:3] != 10'h03E) &&
         (d[12:3] != 10'h03F) &&
         (d[12:3] != 10'h040) &&
         (d[12:3] != 10'h041) &&
         (d[12:3] != 10'h042) &&
         (d[12:3] != 10'h043) &&
         (d[12:3] != 10'h044) &&
         (d[12:3] != 10'h045) &&
         (d[12:3] != 10'h046) &&
         (d[12:3] != 10'h047) &&
         (d[12:3] != 10'h048) &&
         (d[12:3] != 10'h049) &&
         (d[12:3] != 10'h04A) &&
         (d[12:3] != 10'h04B)) ;
  end

initial begin
	$dumpfile( "long_exp2.vcd" );
	$dumpvars( 0, main );
	b = 1'b0;
	c = 1'b0;
	d = 25'h0000000;
	e = 1'b0;
	#5;
	$finish;
end

endmodule

/* HEADER
GROUPS long_exp2 all iv vcs vcd lxt
SIM    long_exp2 all iv vcd  : iverilog long_exp2.v; ./a.out                             : long_exp2.vcd
SIM    long_exp2 all iv lxt  : iverilog long_exp2.v; ./a.out -lxt2; mv long_exp2.vcd long_exp2.lxt : long_exp2.lxt
SIM    long_exp2 all vcs vcd : vcs long_exp2.v; ./simv                                   : long_exp2.vcd
SCORE  long_exp2.vcd     : -t main -vcd long_exp2.vcd -o long_exp2.cdd -v long_exp2.v : long_exp2.cdd
SCORE  long_exp2.lxt     : -t main -lxt long_exp2.lxt -o long_exp2.cdd -v long_exp2.v : long_exp2.cdd
REPORT long_exp2.cdd 1   : -d v -o long_exp2.rptM long_exp2.cdd                         : long_exp2.rptM
REPORT long_exp2.cdd 2   : -d v -w -o long_exp2.rptWM long_exp2.cdd                     : long_exp2.rptWM
REPORT long_exp2.cdd 3   : -d v -i -o long_exp2.rptI long_exp2.cdd                      : long_exp2.rptI
REPORT long_exp2.cdd 4   : -d v -w -i -o long_exp2.rptWI long_exp2.cdd                  : long_exp2.rptWI
*/

/* OUTPUT long_exp2.cdd
5 1 * 6 0 0 0 0
3 0 main main long_exp2.v 1 189
2 1 175 15001b 0 0 20010 0 0 10 3 45 10 0
2 2 175 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 3 175 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 4 175 a0010 0 24 30 2 3 d
2 5 175 a001b 0 15 20030 1 4 1 0 2
2 6 174 15001b 0 0 20010 0 0 10 3 44 10 0
2 7 174 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 8 174 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 9 174 a0010 0 24 30 7 8 d
2 10 174 a001b 0 15 20030 6 9 1 0 2
2 11 173 15001b 0 0 20010 0 0 10 3 41 10 0
2 12 173 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 13 173 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 14 173 a0010 0 24 30 12 13 d
2 15 173 a001b 0 15 20030 11 14 1 0 2
2 16 172 15001b 0 0 20010 0 0 10 3 40 10 0
2 17 172 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 18 172 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 19 172 a0010 0 24 30 17 18 d
2 20 172 a001b 0 15 20030 16 19 1 0 2
2 21 171 15001b 0 0 20010 0 0 10 3 15 10 0
2 22 171 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 23 171 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 24 171 a0010 0 24 30 22 23 d
2 25 171 a001b 0 15 20030 21 24 1 0 2
2 26 170 15001b 0 0 20010 0 0 10 3 14 10 0
2 27 170 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 28 170 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 29 170 a0010 0 24 30 27 28 d
2 30 170 a001b 0 15 20030 26 29 1 0 2
2 31 169 15001b 0 0 20010 0 0 10 3 11 10 0
2 32 169 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 33 169 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 34 169 a0010 0 24 30 32 33 d
2 35 169 a001b 0 15 20030 31 34 1 0 2
2 36 168 15001b 0 0 20010 0 0 10 3 10 10 0
2 37 168 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 38 168 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 39 168 a0010 0 24 30 37 38 d
2 40 168 a001b 0 15 20030 36 39 1 0 2
2 41 167 15001b 0 0 20010 0 0 10 3 5 10 0
2 42 167 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 43 167 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 44 167 a0010 0 24 30 42 43 d
2 45 167 a001b 0 15 20030 41 44 1 0 2
2 46 166 15001b 0 0 20010 0 0 10 3 4 10 0
2 47 166 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 48 166 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 49 166 a0010 0 24 30 47 48 d
2 50 166 a001b 0 15 20030 46 49 1 0 2
2 51 165 15001b 0 0 20010 0 0 10 3 1 10 0
2 52 165 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 53 165 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 54 165 a0010 0 24 30 52 53 d
2 55 165 a001b 0 15 20030 51 54 1 0 2
2 56 164 15001b 0 0 20010 0 0 10 3 0 10 0
2 57 164 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 58 164 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 59 164 a0010 0 24 30 57 58 d
2 60 164 a001b 0 15 20030 56 59 1 0 2
2 61 163 15001b 0 0 20010 0 0 10 3 55 5 0
2 62 163 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 63 163 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 64 163 a0010 0 24 30 62 63 d
2 65 163 a001b 0 15 20030 61 64 1 0 2
2 66 162 15001b 0 0 20010 0 0 10 3 54 5 0
2 67 162 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 68 162 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 69 162 a0010 0 24 30 67 68 d
2 70 162 a001b 0 15 20030 66 69 1 0 2
2 71 161 15001b 0 0 20010 0 0 10 3 51 5 0
2 72 161 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 73 161 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 74 161 a0010 0 24 30 72 73 d
2 75 161 a001b 0 15 20030 71 74 1 0 2
2 76 160 15001b 0 0 20010 0 0 10 3 50 5 0
2 77 160 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 78 160 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 79 160 a0010 0 24 30 77 78 d
2 80 160 a001b 0 15 20030 76 79 1 0 2
2 81 159 15001b 0 0 20010 0 0 10 3 45 5 0
2 82 159 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 83 159 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 84 159 a0010 0 24 30 82 83 d
2 85 159 a001b 0 15 20030 81 84 1 0 2
2 86 158 15001b 0 0 20010 0 0 10 3 44 5 0
2 87 158 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 88 158 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 89 158 a0010 0 24 30 87 88 d
2 90 158 a001b 0 15 20030 86 89 1 0 2
2 91 157 15001b 0 0 20010 0 0 10 3 41 5 0
2 92 157 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 93 157 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 94 157 a0010 0 24 30 92 93 d
2 95 157 a001b 0 15 20030 91 94 1 0 2
2 96 156 15001b 0 0 20010 0 0 10 3 40 5 0
2 97 156 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 98 156 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 99 156 a0010 0 24 30 97 98 d
2 100 156 a001b 0 15 20030 96 99 1 0 2
2 101 155 15001b 0 0 20010 0 0 10 3 15 5 0
2 102 155 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 103 155 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 104 155 a0010 0 24 30 102 103 d
2 105 155 a001b 0 15 20030 101 104 1 0 2
2 106 154 15001b 0 0 20010 0 0 10 3 14 5 0
2 107 154 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 108 154 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 109 154 a0010 0 24 30 107 108 d
2 110 154 a001b 0 15 20030 106 109 1 0 2
2 111 153 15001b 0 0 20010 0 0 10 3 11 5 0
2 112 153 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 113 153 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 114 153 a0010 0 24 30 112 113 d
2 115 153 a001b 0 15 20030 111 114 1 0 2
2 116 152 15001b 0 0 20010 0 0 10 3 10 5 0
2 117 152 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 118 152 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 119 152 a0010 0 24 30 117 118 d
2 120 152 a001b 0 15 20030 116 119 1 0 2
2 121 151 15001b 0 0 20010 0 0 10 3 5 5 0
2 122 151 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 123 151 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 124 151 a0010 0 24 30 122 123 d
2 125 151 a001b 0 15 20030 121 124 1 0 2
2 126 150 15001b 0 0 20010 0 0 10 3 4 5 0
2 127 150 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 128 150 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 129 150 a0010 0 24 30 127 128 d
2 130 150 a001b 0 15 20030 126 129 1 0 2
2 131 149 15001b 0 0 20010 0 0 10 3 1 5 0
2 132 149 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 133 149 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 134 149 a0010 0 24 30 132 133 d
2 135 149 a001b 0 15 20030 131 134 1 0 2
2 136 148 15001b 0 0 20010 0 0 10 3 0 5 0
2 137 148 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 138 148 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 139 148 a0010 0 24 30 137 138 d
2 140 148 a001b 0 15 20030 136 139 1 0 2
2 141 147 15001b 0 0 20010 0 0 10 3 55 4 0
2 142 147 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 143 147 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 144 147 a0010 0 24 30 142 143 d
2 145 147 a001b 0 15 20030 141 144 1 0 2
2 146 146 15001b 0 0 20010 0 0 10 3 54 4 0
2 147 146 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 148 146 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 149 146 a0010 0 24 30 147 148 d
2 150 146 a001b 0 15 20030 146 149 1 0 2
2 151 145 15001b 0 0 20010 0 0 10 3 51 4 0
2 152 145 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 153 145 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 154 145 a0010 0 24 30 152 153 d
2 155 145 a001b 0 15 20030 151 154 1 0 2
2 156 144 15001b 0 0 20010 0 0 10 3 50 4 0
2 157 144 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 158 144 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 159 144 a0010 0 24 30 157 158 d
2 160 144 a001b 0 15 20030 156 159 1 0 2
2 161 143 15001b 0 0 20010 0 0 10 3 45 4 0
2 162 143 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 163 143 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 164 143 a0010 0 24 30 162 163 d
2 165 143 a001b 0 15 20030 161 164 1 0 2
2 166 142 15001b 0 0 20010 0 0 10 3 44 4 0
2 167 142 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 168 142 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 169 142 a0010 0 24 30 167 168 d
2 170 142 a001b 0 15 20030 166 169 1 0 2
2 171 141 15001b 0 0 20010 0 0 10 3 41 4 0
2 172 141 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 173 141 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 174 141 a0010 0 24 30 172 173 d
2 175 141 a001b 0 15 20030 171 174 1 0 2
2 176 140 15001b 0 0 20010 0 0 10 3 40 4 0
2 177 140 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 178 140 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 179 140 a0010 0 24 30 177 178 d
2 180 140 a001b 0 15 20030 176 179 1 0 2
2 181 139 15001b 0 0 20010 0 0 10 3 15 4 0
2 182 139 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 183 139 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 184 139 a0010 0 24 30 182 183 d
2 185 139 a001b 0 15 20030 181 184 1 0 2
2 186 138 15001b 0 0 20010 0 0 10 3 14 4 0
2 187 138 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 188 138 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 189 138 a0010 0 24 30 187 188 d
2 190 138 a001b 0 15 20030 186 189 1 0 2
2 191 137 15001b 0 0 20010 0 0 10 3 11 4 0
2 192 137 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 193 137 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 194 137 a0010 0 24 30 192 193 d
2 195 137 a001b 0 15 20030 191 194 1 0 2
2 196 136 15001b 0 0 20010 0 0 10 3 10 4 0
2 197 136 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 198 136 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 199 136 a0010 0 24 30 197 198 d
2 200 136 a001b 0 15 20030 196 199 1 0 2
2 201 135 15001b 0 0 20010 0 0 10 3 5 4 0
2 202 135 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 203 135 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 204 135 a0010 0 24 30 202 203 d
2 205 135 a001b 0 15 20030 201 204 1 0 2
2 206 134 15001b 0 0 20010 0 0 10 3 4 4 0
2 207 134 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 208 134 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 209 134 a0010 0 24 30 207 208 d
2 210 134 a001b 0 15 20030 206 209 1 0 2
2 211 133 15001b 0 0 20010 0 0 10 3 1 4 0
2 212 133 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 213 133 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 214 133 a0010 0 24 30 212 213 d
2 215 133 a001b 0 15 20030 211 214 1 0 2
2 216 132 15001b 0 0 20010 0 0 10 3 0 4 0
2 217 132 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 218 132 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 219 132 a0010 0 24 30 217 218 d
2 220 132 a001b 0 15 20030 216 219 1 0 2
2 221 131 15001b 0 0 20010 0 0 10 3 55 1 0
2 222 131 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 223 131 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 224 131 a0010 0 24 30 222 223 d
2 225 131 a001b 0 15 20030 221 224 1 0 2
2 226 130 15001b 0 0 20010 0 0 10 3 54 1 0
2 227 130 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 228 130 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 229 130 a0010 0 24 30 227 228 d
2 230 130 a001b 0 15 20030 226 229 1 0 2
2 231 129 15001b 0 0 20010 0 0 10 3 51 1 0
2 232 129 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 233 129 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 234 129 a0010 0 24 30 232 233 d
2 235 129 a001b 0 15 20030 231 234 1 0 2
2 236 128 15001b 0 0 20010 0 0 10 3 50 1 0
2 237 128 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 238 128 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 239 128 a0010 0 24 30 237 238 d
2 240 128 a001b 0 15 20030 236 239 1 0 2
2 241 127 15001b 0 0 20010 0 0 10 3 45 1 0
2 242 127 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 243 127 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 244 127 a0010 0 24 30 242 243 d
2 245 127 a001b 0 15 20030 241 244 1 0 2
2 246 126 15001b 0 0 20010 0 0 10 3 44 1 0
2 247 126 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 248 126 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 249 126 a0010 0 24 30 247 248 d
2 250 126 a001b 0 15 20030 246 249 1 0 2
2 251 125 15001b 0 0 20010 0 0 10 3 41 1 0
2 252 125 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 253 125 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 254 125 a0010 0 24 30 252 253 d
2 255 125 a001b 0 15 20030 251 254 1 0 2
2 256 124 15001b 0 0 20010 0 0 10 3 40 1 0
2 257 124 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 258 124 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 259 124 a0010 0 24 30 257 258 d
2 260 124 a001b 0 15 20030 256 259 1 0 2
2 261 123 15001b 0 0 20010 0 0 10 3 15 1 0
2 262 123 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 263 123 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 264 123 a0010 0 24 30 262 263 d
2 265 123 a001b 0 15 20030 261 264 1 0 2
2 266 122 15001b 0 0 20010 0 0 10 3 14 1 0
2 267 122 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 268 122 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 269 122 a0010 0 24 30 267 268 d
2 270 122 a001b 0 15 20030 266 269 1 0 2
2 271 121 15001b 0 0 20010 0 0 10 3 11 1 0
2 272 121 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 273 121 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 274 121 a0010 0 24 30 272 273 d
2 275 121 a001b 0 15 20030 271 274 1 0 2
2 276 120 15001b 0 0 20010 0 0 10 3 10 1 0
2 277 120 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 278 120 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 279 120 a0010 0 24 30 277 278 d
2 280 120 a001b 0 15 20030 276 279 1 0 2
2 281 119 15001b 0 0 20010 0 0 10 3 5 1 0
2 282 119 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 283 119 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 284 119 a0010 0 24 30 282 283 d
2 285 119 a001b 0 15 20030 281 284 1 0 2
2 286 118 15001b 0 0 20010 0 0 10 3 4 1 0
2 287 118 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 288 118 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 289 118 a0010 0 24 30 287 288 d
2 290 118 a001b 0 15 20030 286 289 1 0 2
2 291 117 15001b 0 0 20010 0 0 10 3 1 1 0
2 292 117 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 293 117 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 294 117 a0010 0 24 30 292 293 d
2 295 117 a001b 0 15 20030 291 294 1 0 2
2 296 116 15001b 0 0 20010 0 0 10 3 0 1 0
2 297 116 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 298 116 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 299 116 a0010 0 24 30 297 298 d
2 300 116 a001b 0 15 20030 296 299 1 0 2
2 301 115 15001b 0 0 20010 0 0 10 3 55 0 0
2 302 115 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 303 115 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 304 115 a0010 0 24 30 302 303 d
2 305 115 a001b 0 15 20030 301 304 1 0 2
2 306 114 15001b 0 0 20010 0 0 10 3 54 0 0
2 307 114 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 308 114 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 309 114 a0010 0 24 30 307 308 d
2 310 114 a001b 0 15 20030 306 309 1 0 2
2 311 113 15001b 0 0 20010 0 0 10 3 51 0 0
2 312 113 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 313 113 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 314 113 a0010 0 24 30 312 313 d
2 315 113 a001b 0 15 20030 311 314 1 0 2
2 316 112 15001b 0 0 20010 0 0 10 3 50 0 0
2 317 112 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 318 112 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 319 112 a0010 0 24 30 317 318 d
2 320 112 a001b 0 15 20030 316 319 1 0 2
2 321 111 15001b 0 0 20010 0 0 10 3 45 0 0
2 322 111 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 323 111 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 324 111 a0010 0 24 30 322 323 d
2 325 111 a001b 0 15 20030 321 324 1 0 2
2 326 110 15001b 0 0 20010 0 0 10 3 44 0 0
2 327 110 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 328 110 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 329 110 a0010 0 24 30 327 328 d
2 330 110 a001b 0 15 20030 326 329 1 0 2
2 331 109 15001b 0 0 20010 0 0 10 3 41 0 0
2 332 109 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 333 109 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 334 109 a0010 0 24 30 332 333 d
2 335 109 a001b 0 15 20030 331 334 1 0 2
2 336 108 15001b 0 0 20010 0 0 10 3 40 0 0
2 337 108 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 338 108 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 339 108 a0010 0 24 30 337 338 d
2 340 108 a001b 0 15 20030 336 339 1 0 2
2 341 107 15001b 0 0 20010 0 0 10 3 15 0 0
2 342 107 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 343 107 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 344 107 a0010 0 24 30 342 343 d
2 345 107 a001b 0 15 20030 341 344 1 0 2
2 346 106 15001b 0 0 20010 0 0 10 3 14 0 0
2 347 106 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 348 106 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 349 106 a0010 0 24 30 347 348 d
2 350 106 a001b 0 15 20030 346 349 1 0 2
2 351 105 15001b 0 0 20010 0 0 10 3 11 0 0
2 352 105 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 353 105 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 354 105 a0010 0 24 30 352 353 d
2 355 105 a001b 0 15 20030 351 354 1 0 2
2 356 104 15001b 0 0 20010 0 0 10 3 10 0 0
2 357 104 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 358 104 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 359 104 a0010 0 24 30 357 358 d
2 360 104 a001b 0 15 20030 356 359 1 0 2
2 361 103 15001b 0 0 20010 0 0 10 3 5 0 0
2 362 103 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 363 103 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 364 103 a0010 0 24 30 362 363 d
2 365 103 a001b 0 15 20030 361 364 1 0 2
2 366 102 15001b 0 0 20010 0 0 10 3 4 0 0
2 367 102 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 368 102 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 369 102 a0010 0 24 30 367 368 d
2 370 102 a001b 0 15 20030 366 369 1 0 2
2 371 101 15001b 0 0 20010 0 0 10 3 1 0 0
2 372 101 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 373 101 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 374 101 a0010 0 24 30 372 373 d
2 375 101 a001b 0 15 20030 371 374 1 0 2
2 376 100 15001b 0 0 20010 0 0 10 3 0 0 0
2 377 100 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 378 100 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 379 100 a0010 0 24 30 377 378 d
2 380 100 a001b 0 15 20030 376 379 1 0 2
2 381 99 140018 0 0 20010 0 0 12 3 0 0 0
2 382 99 f0010 0 0 20018 0 0 32 64 0 1 0 0 0 0 0 0
2 383 99 c000d 0 0 20018 0 0 32 64 45 1 0 0 0 0 0 0
2 384 99 a0011 0 24 30 382 383 d
2 385 99 a0018 0 11 20030 381 384 1 0 2
2 386 99 9001c 0 18 20030 380 385 1 0 2
2 387 99 9001c 0 18 20030 375 386 1 0 2
2 388 99 9001c 0 18 20030 370 387 1 0 2
2 389 99 9001c 0 18 20030 365 388 1 0 2
2 390 99 9001c 0 18 20030 360 389 1 0 2
2 391 99 9001c 0 18 20030 355 390 1 0 2
2 392 99 9001c 0 18 20030 350 391 1 0 2
2 393 99 9001c 0 18 20030 345 392 1 0 2
2 394 99 9001c 0 18 20030 340 393 1 0 2
2 395 99 9001c 0 18 20030 335 394 1 0 2
2 396 99 9001c 0 18 20030 330 395 1 0 2
2 397 99 9001c 0 18 20030 325 396 1 0 2
2 398 99 9001c 0 18 20030 320 397 1 0 2
2 399 99 9001c 0 18 20030 315 398 1 0 2
2 400 99 9001c 0 18 20030 310 399 1 0 2
2 401 99 9001c 0 18 20030 305 400 1 0 2
2 402 99 9001c 0 18 20030 300 401 1 0 2
2 403 99 9001c 0 18 20030 295 402 1 0 2
2 404 99 9001c 0 18 20030 290 403 1 0 2
2 405 99 9001c 0 18 20030 285 404 1 0 2
2 406 99 9001c 0 18 20030 280 405 1 0 2
2 407 99 9001c 0 18 20030 275 406 1 0 2
2 408 99 9001c 0 18 20030 270 407 1 0 2
2 409 99 9001c 0 18 20030 265 408 1 0 2
2 410 99 9001c 0 18 20030 260 409 1 0 2
2 411 99 9001c 0 18 20030 255 410 1 0 2
2 412 99 9001c 0 18 20030 250 411 1 0 2
2 413 99 9001c 0 18 20030 245 412 1 0 2
2 414 99 9001c 0 18 20030 240 413 1 0 2
2 415 99 9001c 0 18 20030 235 414 1 0 2
2 416 99 9001c 0 18 20030 230 415 1 0 2
2 417 99 9001c 0 18 20030 225 416 1 0 2
2 418 99 9001c 0 18 20030 220 417 1 0 2
2 419 99 9001c 0 18 20030 215 418 1 0 2
2 420 99 9001c 0 18 20030 210 419 1 0 2
2 421 99 9001c 0 18 20030 205 420 1 0 2
2 422 99 9001c 0 18 20030 200 421 1 0 2
2 423 99 9001c 0 18 20030 195 422 1 0 2
2 424 99 9001c 0 18 20030 190 423 1 0 2
2 425 99 9001c 0 18 20030 185 424 1 0 2
2 426 99 9001c 0 18 20030 180 425 1 0 2
2 427 99 9001c 0 18 20030 175 426 1 0 2
2 428 99 9001c 0 18 20030 170 427 1 0 2
2 429 99 9001c 0 18 20030 165 428 1 0 2
2 430 99 9001c 0 18 20030 160 429 1 0 2
2 431 99 9001c 0 18 20030 155 430 1 0 2
2 432 99 9001c 0 18 20030 150 431 1 0 2
2 433 99 9001c 0 18 20030 145 432 1 0 2
2 434 99 9001c 0 18 20030 140 433 1 0 2
2 435 99 9001c 0 18 20030 135 434 1 0 2
2 436 99 9001c 0 18 20030 130 435 1 0 2
2 437 99 9001c 0 18 20030 125 436 1 0 2
2 438 99 9001c 0 18 20030 120 437 1 0 2
2 439 99 9001c 0 18 20030 115 438 1 0 2
2 440 99 9001c 0 18 20030 110 439 1 0 2
2 441 99 9001c 0 18 20030 105 440 1 0 2
2 442 99 9001c 0 18 20030 100 441 1 0 2
2 443 99 9001c 0 18 20030 95 442 1 0 2
2 444 99 9001c 0 18 20030 90 443 1 0 2
2 445 99 9001c 0 18 20030 85 444 1 0 2
2 446 99 9001c 0 18 20030 80 445 1 0 2
2 447 99 9001c 0 18 20030 75 446 1 0 2
2 448 99 9001c 0 18 20030 70 447 1 0 2
2 449 99 9001c 0 18 20030 65 448 1 0 2
2 450 99 9001c 0 18 20030 60 449 1 0 2
2 451 99 9001c 0 18 20030 55 450 1 0 2
2 452 99 9001c 0 18 20030 50 451 1 0 2
2 453 99 9001c 0 18 20030 45 452 1 0 2
2 454 99 9001c 0 18 20030 40 453 1 0 2
2 455 99 9001c 0 18 20030 35 454 1 0 2
2 456 99 9001c 0 18 20030 30 455 1 0 2
2 457 99 9001c 0 18 20030 25 456 1 0 2
2 458 99 9001c 0 18 20030 20 457 1 0 2
2 459 99 9001c 0 18 20030 15 458 1 0 2
2 460 99 9001c 0 18 20030 10 459 1 0 2
2 461 99 9001c 0 18 20030 5 460 1 0 2
2 462 98 80008 0 1 10 0 0 e
2 463 98 8001d 0 8 20030 461 462 1 0 2
2 464 97 15001b 0 0 20010 0 0 10 3 10 11 0
2 465 97 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 466 97 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 467 97 a0010 0 24 30 465 466 d
2 468 97 a001b 0 15 20030 464 467 1 0 2
2 469 96 15001b 0 0 20010 0 0 10 3 5 11 0
2 470 96 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 471 96 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 472 96 a0010 0 24 30 470 471 d
2 473 96 a001b 0 15 20030 469 472 1 0 2
2 474 95 15001b 0 0 20010 0 0 10 3 4 11 0
2 475 95 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 476 95 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 477 95 a0010 0 24 30 475 476 d
2 478 95 a001b 0 15 20030 474 477 1 0 2
2 479 94 15001b 0 0 20010 0 0 10 3 1 11 0
2 480 94 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 481 94 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 482 94 a0010 0 24 30 480 481 d
2 483 94 a001b 0 15 20030 479 482 1 0 2
2 484 93 15001b 0 0 20010 0 0 10 3 0 11 0
2 485 93 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 486 93 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 487 93 a0010 0 24 30 485 486 d
2 488 93 a001b 0 15 20030 484 487 1 0 2
2 489 92 15001b 0 0 20010 0 0 10 3 55 10 0
2 490 92 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 491 92 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 492 92 a0010 0 24 30 490 491 d
2 493 92 a001b 0 15 20030 489 492 1 0 2
2 494 91 15001b 0 0 20010 0 0 10 3 54 10 0
2 495 91 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 496 91 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 497 91 a0010 0 24 30 495 496 d
2 498 91 a001b 0 15 20030 494 497 1 0 2
2 499 90 15001b 0 0 20010 0 0 10 3 51 10 0
2 500 90 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 501 90 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 502 90 a0010 0 24 30 500 501 d
2 503 90 a001b 0 15 20030 499 502 1 0 2
2 504 89 15001b 0 0 20010 0 0 10 3 50 10 0
2 505 89 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 506 89 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 507 89 a0010 0 24 30 505 506 d
2 508 89 a001b 0 15 20030 504 507 1 0 2
2 509 88 15001b 0 0 20010 0 0 10 3 45 10 0
2 510 88 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 511 88 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 512 88 a0010 0 24 30 510 511 d
2 513 88 a001b 0 15 20030 509 512 1 0 2
2 514 87 15001b 0 0 20010 0 0 10 3 44 10 0
2 515 87 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 516 87 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 517 87 a0010 0 24 30 515 516 d
2 518 87 a001b 0 15 20030 514 517 1 0 2
2 519 86 15001b 0 0 20010 0 0 10 3 41 10 0
2 520 86 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 521 86 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 522 86 a0010 0 24 30 520 521 d
2 523 86 a001b 0 15 20030 519 522 1 0 2
2 524 85 15001b 0 0 20010 0 0 10 3 40 10 0
2 525 85 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 526 85 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 527 85 a0010 0 24 30 525 526 d
2 528 85 a001b 0 15 20030 524 527 1 0 2
2 529 84 15001b 0 0 20010 0 0 10 3 15 10 0
2 530 84 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 531 84 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 532 84 a0010 0 24 30 530 531 d
2 533 84 a001b 0 15 20030 529 532 1 0 2
2 534 83 15001b 0 0 20010 0 0 10 3 14 10 0
2 535 83 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 536 83 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 537 83 a0010 0 24 30 535 536 d
2 538 83 a001b 0 15 20030 534 537 1 0 2
2 539 82 15001b 0 0 20010 0 0 10 3 11 10 0
2 540 82 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 541 82 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 542 82 a0010 0 24 30 540 541 d
2 543 82 a001b 0 15 20030 539 542 1 0 2
2 544 81 15001b 0 0 20010 0 0 10 3 10 10 0
2 545 81 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 546 81 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 547 81 a0010 0 24 30 545 546 d
2 548 81 a001b 0 15 20030 544 547 1 0 2
2 549 80 15001b 0 0 20010 0 0 10 3 5 10 0
2 550 80 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 551 80 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 552 80 a0010 0 24 30 550 551 d
2 553 80 a001b 0 15 20030 549 552 1 0 2
2 554 79 15001b 0 0 20010 0 0 10 3 4 10 0
2 555 79 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 556 79 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 557 79 a0010 0 24 30 555 556 d
2 558 79 a001b 0 15 20030 554 557 1 0 2
2 559 78 15001b 0 0 20010 0 0 10 3 1 10 0
2 560 78 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 561 78 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 562 78 a0010 0 24 30 560 561 d
2 563 78 a001b 0 15 20030 559 562 1 0 2
2 564 77 15001b 0 0 20010 0 0 10 3 0 10 0
2 565 77 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 566 77 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 567 77 a0010 0 24 30 565 566 d
2 568 77 a001b 0 15 20030 564 567 1 0 2
2 569 76 15001b 0 0 20010 0 0 10 3 55 5 0
2 570 76 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 571 76 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 572 76 a0010 0 24 30 570 571 d
2 573 76 a001b 0 15 20030 569 572 1 0 2
2 574 75 15001b 0 0 20010 0 0 10 3 54 5 0
2 575 75 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 576 75 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 577 75 a0010 0 24 30 575 576 d
2 578 75 a001b 0 15 20030 574 577 1 0 2
2 579 74 15001b 0 0 20010 0 0 10 3 51 5 0
2 580 74 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 581 74 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 582 74 a0010 0 24 30 580 581 d
2 583 74 a001b 0 15 20030 579 582 1 0 2
2 584 73 15001b 0 0 20010 0 0 10 3 50 5 0
2 585 73 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 586 73 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 587 73 a0010 0 24 30 585 586 d
2 588 73 a001b 0 15 20030 584 587 1 0 2
2 589 72 15001b 0 0 20010 0 0 10 3 45 5 0
2 590 72 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 591 72 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 592 72 a0010 0 24 30 590 591 d
2 593 72 a001b 0 15 20030 589 592 1 0 2
2 594 71 15001b 0 0 20010 0 0 10 3 44 5 0
2 595 71 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 596 71 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 597 71 a0010 0 24 30 595 596 d
2 598 71 a001b 0 15 20030 594 597 1 0 2
2 599 70 15001b 0 0 20010 0 0 10 3 41 5 0
2 600 70 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 601 70 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 602 70 a0010 0 24 30 600 601 d
2 603 70 a001b 0 15 20030 599 602 1 0 2
2 604 69 15001b 0 0 20010 0 0 10 3 40 5 0
2 605 69 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 606 69 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 607 69 a0010 0 24 30 605 606 d
2 608 69 a001b 0 15 20030 604 607 1 0 2
2 609 68 15001b 0 0 20010 0 0 10 3 15 5 0
2 610 68 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 611 68 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 612 68 a0010 0 24 30 610 611 d
2 613 68 a001b 0 15 20030 609 612 1 0 2
2 614 67 15001b 0 0 20010 0 0 10 3 14 5 0
2 615 67 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 616 67 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 617 67 a0010 0 24 30 615 616 d
2 618 67 a001b 0 15 20030 614 617 1 0 2
2 619 66 15001b 0 0 20010 0 0 10 3 11 5 0
2 620 66 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 621 66 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 622 66 a0010 0 24 30 620 621 d
2 623 66 a001b 0 15 20030 619 622 1 0 2
2 624 65 15001b 0 0 20010 0 0 10 3 10 5 0
2 625 65 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 626 65 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 627 65 a0010 0 24 30 625 626 d
2 628 65 a001b 0 15 20030 624 627 1 0 2
2 629 64 15001b 0 0 20010 0 0 10 3 5 5 0
2 630 64 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 631 64 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 632 64 a0010 0 24 30 630 631 d
2 633 64 a001b 0 15 20030 629 632 1 0 2
2 634 63 15001b 0 0 20010 0 0 10 3 4 5 0
2 635 63 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 636 63 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 637 63 a0010 0 24 30 635 636 d
2 638 63 a001b 0 15 20030 634 637 1 0 2
2 639 62 15001b 0 0 20010 0 0 10 3 1 5 0
2 640 62 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 641 62 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 642 62 a0010 0 24 30 640 641 d
2 643 62 a001b 0 15 20030 639 642 1 0 2
2 644 61 15001b 0 0 20010 0 0 10 3 0 5 0
2 645 61 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 646 61 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 647 61 a0010 0 24 30 645 646 d
2 648 61 a001b 0 15 20030 644 647 1 0 2
2 649 60 15001b 0 0 20010 0 0 10 3 55 4 0
2 650 60 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 651 60 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 652 60 a0010 0 24 30 650 651 d
2 653 60 a001b 0 15 20030 649 652 1 0 2
2 654 59 15001b 0 0 20010 0 0 10 3 54 4 0
2 655 59 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 656 59 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 657 59 a0010 0 24 30 655 656 d
2 658 59 a001b 0 15 20030 654 657 1 0 2
2 659 58 15001b 0 0 20010 0 0 10 3 51 4 0
2 660 58 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 661 58 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 662 58 a0010 0 24 30 660 661 d
2 663 58 a001b 0 15 20030 659 662 1 0 2
2 664 57 15001b 0 0 20010 0 0 10 3 50 4 0
2 665 57 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 666 57 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 667 57 a0010 0 24 30 665 666 d
2 668 57 a001b 0 15 20030 664 667 1 0 2
2 669 56 15001b 0 0 20010 0 0 10 3 45 4 0
2 670 56 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 671 56 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 672 56 a0010 0 24 30 670 671 d
2 673 56 a001b 0 15 20030 669 672 1 0 2
2 674 55 15001b 0 0 20010 0 0 10 3 44 4 0
2 675 55 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 676 55 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 677 55 a0010 0 24 30 675 676 d
2 678 55 a001b 0 15 20030 674 677 1 0 2
2 679 54 15001b 0 0 20010 0 0 10 3 41 4 0
2 680 54 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 681 54 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 682 54 a0010 0 24 30 680 681 d
2 683 54 a001b 0 15 20030 679 682 1 0 2
2 684 53 15001b 0 0 20010 0 0 10 3 40 4 0
2 685 53 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 686 53 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 687 53 a0010 0 24 30 685 686 d
2 688 53 a001b 0 15 20030 684 687 1 0 2
2 689 52 15001b 0 0 20010 0 0 10 3 15 4 0
2 690 52 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 691 52 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 692 52 a0010 0 24 30 690 691 d
2 693 52 a001b 0 15 20030 689 692 1 0 2
2 694 51 15001b 0 0 20010 0 0 10 3 14 4 0
2 695 51 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 696 51 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 697 51 a0010 0 24 30 695 696 d
2 698 51 a001b 0 15 20030 694 697 1 0 2
2 699 50 15001b 0 0 20010 0 0 10 3 11 4 0
2 700 50 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 701 50 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 702 50 a0010 0 24 30 700 701 d
2 703 50 a001b 0 15 20030 699 702 1 0 2
2 704 49 15001b 0 0 20010 0 0 10 3 10 4 0
2 705 49 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 706 49 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 707 49 a0010 0 24 30 705 706 d
2 708 49 a001b 0 15 20030 704 707 1 0 2
2 709 48 15001b 0 0 20010 0 0 10 3 5 4 0
2 710 48 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 711 48 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 712 48 a0010 0 24 30 710 711 d
2 713 48 a001b 0 15 20030 709 712 1 0 2
2 714 47 15001b 0 0 20010 0 0 10 3 4 4 0
2 715 47 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 716 47 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 717 47 a0010 0 24 30 715 716 d
2 718 47 a001b 0 15 20030 714 717 1 0 2
2 719 46 15001b 0 0 20010 0 0 10 3 1 4 0
2 720 46 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 721 46 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 722 46 a0010 0 24 30 720 721 d
2 723 46 a001b 0 15 20030 719 722 1 0 2
2 724 45 15001b 0 0 20010 0 0 10 3 0 4 0
2 725 45 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 726 45 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 727 45 a0010 0 24 30 725 726 d
2 728 45 a001b 0 15 20030 724 727 1 0 2
2 729 44 15001b 0 0 20010 0 0 10 3 55 1 0
2 730 44 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 731 44 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 732 44 a0010 0 24 30 730 731 d
2 733 44 a001b 0 15 20030 729 732 1 0 2
2 734 43 15001b 0 0 20010 0 0 10 3 54 1 0
2 735 43 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 736 43 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 737 43 a0010 0 24 30 735 736 d
2 738 43 a001b 0 15 20030 734 737 1 0 2
2 739 42 15001b 0 0 20010 0 0 10 3 51 1 0
2 740 42 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 741 42 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 742 42 a0010 0 24 30 740 741 d
2 743 42 a001b 0 15 20030 739 742 1 0 2
2 744 41 15001b 0 0 20010 0 0 10 3 50 1 0
2 745 41 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 746 41 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 747 41 a0010 0 24 30 745 746 d
2 748 41 a001b 0 15 20030 744 747 1 0 2
2 749 40 15001b 0 0 20010 0 0 10 3 45 1 0
2 750 40 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 751 40 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 752 40 a0010 0 24 30 750 751 d
2 753 40 a001b 0 15 20030 749 752 1 0 2
2 754 39 15001b 0 0 20010 0 0 10 3 44 1 0
2 755 39 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 756 39 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 757 39 a0010 0 24 30 755 756 d
2 758 39 a001b 0 15 20030 754 757 1 0 2
2 759 38 15001b 0 0 20010 0 0 10 3 41 1 0
2 760 38 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 761 38 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 762 38 a0010 0 24 30 760 761 d
2 763 38 a001b 0 15 20030 759 762 1 0 2
2 764 37 15001b 0 0 20010 0 0 10 3 40 1 0
2 765 37 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 766 37 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 767 37 a0010 0 24 30 765 766 d
2 768 37 a001b 0 15 20030 764 767 1 0 2
2 769 36 15001b 0 0 20010 0 0 10 3 15 1 0
2 770 36 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 771 36 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 772 36 a0010 0 24 30 770 771 d
2 773 36 a001b 0 15 20030 769 772 1 0 2
2 774 35 15001b 0 0 20010 0 0 10 3 14 1 0
2 775 35 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 776 35 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 777 35 a0010 0 24 30 775 776 d
2 778 35 a001b 0 15 20030 774 777 1 0 2
2 779 34 15001b 0 0 20010 0 0 10 3 11 1 0
2 780 34 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 781 34 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 782 34 a0010 0 24 30 780 781 d
2 783 34 a001b 0 15 20030 779 782 1 0 2
2 784 33 15001b 0 0 20010 0 0 10 3 10 1 0
2 785 33 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 786 33 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 787 33 a0010 0 24 30 785 786 d
2 788 33 a001b 0 15 20030 784 787 1 0 2
2 789 32 15001b 0 0 20010 0 0 10 3 5 1 0
2 790 32 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 791 32 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 792 32 a0010 0 24 30 790 791 d
2 793 32 a001b 0 15 20030 789 792 1 0 2
2 794 31 15001b 0 0 20010 0 0 10 3 4 1 0
2 795 31 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 796 31 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 797 31 a0010 0 24 30 795 796 d
2 798 31 a001b 0 15 20030 794 797 1 0 2
2 799 30 15001b 0 0 20010 0 0 10 3 1 1 0
2 800 30 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 801 30 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 802 30 a0010 0 24 30 800 801 d
2 803 30 a001b 0 15 20030 799 802 1 0 2
2 804 29 15001b 0 0 20010 0 0 10 3 0 1 0
2 805 29 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 806 29 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 807 29 a0010 0 24 30 805 806 d
2 808 29 a001b 0 15 20030 804 807 1 0 2
2 809 28 15001b 0 0 20010 0 0 10 3 55 0 0
2 810 28 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 811 28 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 812 28 a0010 0 24 30 810 811 d
2 813 28 a001b 0 15 20030 809 812 1 0 2
2 814 27 15001b 0 0 20010 0 0 10 3 54 0 0
2 815 27 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 816 27 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 817 27 a0010 0 24 30 815 816 d
2 818 27 a001b 0 15 20030 814 817 1 0 2
2 819 26 15001b 0 0 20010 0 0 10 3 51 0 0
2 820 26 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 821 26 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 822 26 a0010 0 24 30 820 821 d
2 823 26 a001b 0 15 20030 819 822 1 0 2
2 824 25 15001b 0 0 20010 0 0 10 3 50 0 0
2 825 25 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 826 25 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 827 25 a0010 0 24 30 825 826 d
2 828 25 a001b 0 15 20030 824 827 1 0 2
2 829 24 15001b 0 0 20010 0 0 10 3 45 0 0
2 830 24 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 831 24 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 832 24 a0010 0 24 30 830 831 d
2 833 24 a001b 0 15 20030 829 832 1 0 2
2 834 23 15001b 0 0 20010 0 0 10 3 44 0 0
2 835 23 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 836 23 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 837 23 a0010 0 24 30 835 836 d
2 838 23 a001b 0 15 20030 834 837 1 0 2
2 839 22 15001b 0 0 20010 0 0 10 3 41 0 0
2 840 22 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 841 22 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 842 22 a0010 0 24 30 840 841 d
2 843 22 a001b 0 15 20030 839 842 1 0 2
2 844 21 15001b 0 0 20010 0 0 10 3 40 0 0
2 845 21 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 846 21 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 847 21 a0010 0 24 30 845 846 d
2 848 21 a001b 0 15 20030 844 847 1 0 2
2 849 20 15001b 0 0 20010 0 0 10 3 15 0 0
2 850 20 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 851 20 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 852 20 a0010 0 24 30 850 851 d
2 853 20 a001b 0 15 20030 849 852 1 0 2
2 854 19 15001b 0 0 20010 0 0 10 3 14 0 0
2 855 19 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 856 19 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 857 19 a0010 0 24 30 855 856 d
2 858 19 a001b 0 15 20030 854 857 1 0 2
2 859 18 15001b 0 0 20010 0 0 10 3 11 0 0
2 860 18 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 861 18 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 862 18 a0010 0 24 30 860 861 d
2 863 18 a001b 0 15 20030 859 862 1 0 2
2 864 17 15001b 0 0 20010 0 0 10 3 10 0 0
2 865 17 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 866 17 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 867 17 a0010 0 24 30 865 866 d
2 868 17 a001b 0 15 20030 864 867 1 0 2
2 869 16 15001b 0 0 20010 0 0 10 3 5 0 0
2 870 16 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 871 16 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 872 16 a0010 0 24 30 870 871 d
2 873 16 a001b 0 15 20030 869 872 1 0 2
2 874 15 15001b 0 0 20010 0 0 10 3 4 0 0
2 875 15 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 876 15 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 877 15 a0010 0 24 30 875 876 d
2 878 15 a001b 0 15 20030 874 877 1 0 2
2 879 14 15001b 0 0 20010 0 0 10 3 1 0 0
2 880 14 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 881 14 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 882 14 a0010 0 24 30 880 881 d
2 883 14 a001b 0 15 20030 879 882 1 0 2
2 884 13 15001b 0 0 20010 0 0 10 3 0 0 0
2 885 13 f000f 0 0 20018 0 0 32 64 5 0 0 0 0 0 0 0
2 886 13 c000d 0 0 20018 0 0 32 64 50 0 0 0 0 0 0 0
2 887 13 a0010 0 24 30 885 886 d
2 888 13 a001b 0 15 20030 884 887 1 0 2
2 889 12 150019 0 0 20010 0 0 12 3 0 0 0
2 890 12 100011 0 0 20018 0 0 32 64 0 1 0 0 0 0 0 0
2 891 12 d000e 0 0 20018 0 0 32 64 45 1 0 0 0 0 0 0
2 892 12 b0012 0 24 30 890 891 d
2 893 12 b0019 0 11 20030 889 892 1 0 2
2 894 12 a001c 0 18 20030 888 893 1 0 2
2 895 12 a001c 0 18 20030 883 894 1 0 2
2 896 12 a001c 0 18 20030 878 895 1 0 2
2 897 12 a001c 0 18 20030 873 896 1 0 2
2 898 12 a001c 0 18 20030 868 897 1 0 2
2 899 12 a001c 0 18 20030 863 898 1 0 2
2 900 12 a001c 0 18 20030 858 899 1 0 2
2 901 12 a001c 0 18 20030 853 900 1 0 2
2 902 12 a001c 0 18 20030 848 901 1 0 2
2 903 12 a001c 0 18 20030 843 902 1 0 2
2 904 12 a001c 0 18 20030 838 903 1 0 2
2 905 12 a001c 0 18 20030 833 904 1 0 2
2 906 12 a001c 0 18 20030 828 905 1 0 2
2 907 12 a001c 0 18 20030 823 906 1 0 2
2 908 12 a001c 0 18 20030 818 907 1 0 2
2 909 12 a001c 0 18 20030 813 908 1 0 2
2 910 12 a001c 0 18 20030 808 909 1 0 2
2 911 12 a001c 0 18 20030 803 910 1 0 2
2 912 12 a001c 0 18 20030 798 911 1 0 2
2 913 12 a001c 0 18 20030 793 912 1 0 2
2 914 12 a001c 0 18 20030 788 913 1 0 2
2 915 12 a001c 0 18 20030 783 914 1 0 2
2 916 12 a001c 0 18 20030 778 915 1 0 2
2 917 12 a001c 0 18 20030 773 916 1 0 2
2 918 12 a001c 0 18 20030 768 917 1 0 2
2 919 12 a001c 0 18 20030 763 918 1 0 2
2 920 12 a001c 0 18 20030 758 919 1 0 2
2 921 12 a001c 0 18 20030 753 920 1 0 2
2 922 12 a001c 0 18 20030 748 921 1 0 2
2 923 12 a001c 0 18 20030 743 922 1 0 2
2 924 12 a001c 0 18 20030 738 923 1 0 2
2 925 12 a001c 0 18 20030 733 924 1 0 2
2 926 12 a001c 0 18 20030 728 925 1 0 2
2 927 12 a001c 0 18 20030 723 926 1 0 2
2 928 12 a001c 0 18 20030 718 927 1 0 2
2 929 12 a001c 0 18 20030 713 928 1 0 2
2 930 12 a001c 0 18 20030 708 929 1 0 2
2 931 12 a001c 0 18 20030 703 930 1 0 2
2 932 12 a001c 0 18 20030 698 931 1 0 2
2 933 12 a001c 0 18 20030 693 932 1 0 2
2 934 12 a001c 0 18 20030 688 933 1 0 2
2 935 12 a001c 0 18 20030 683 934 1 0 2
2 936 12 a001c 0 18 20030 678 935 1 0 2
2 937 12 a001c 0 18 20030 673 936 1 0 2
2 938 12 a001c 0 18 20030 668 937 1 0 2
2 939 12 a001c 0 18 20030 663 938 1 0 2
2 940 12 a001c 0 18 20030 658 939 1 0 2
2 941 12 a001c 0 18 20030 653 940 1 0 2
2 942 12 a001c 0 18 20030 648 941 1 0 2
2 943 12 a001c 0 18 20030 643 942 1 0 2
2 944 12 a001c 0 18 20030 638 943 1 0 2
2 945 12 a001c 0 18 20030 633 944 1 0 2
2 946 12 a001c 0 18 20030 628 945 1 0 2
2 947 12 a001c 0 18 20030 623 946 1 0 2
2 948 12 a001c 0 18 20030 618 947 1 0 2
2 949 12 a001c 0 18 20030 613 948 1 0 2
2 950 12 a001c 0 18 20030 608 949 1 0 2
2 951 12 a001c 0 18 20030 603 950 1 0 2
2 952 12 a001c 0 18 20030 598 951 1 0 2
2 953 12 a001c 0 18 20030 593 952 1 0 2
2 954 12 a001c 0 18 20030 588 953 1 0 2
2 955 12 a001c 0 18 20030 583 954 1 0 2
2 956 12 a001c 0 18 20030 578 955 1 0 2
2 957 12 a001c 0 18 20030 573 956 1 0 2
2 958 12 a001c 0 18 20030 568 957 1 0 2
2 959 12 a001c 0 18 20030 563 958 1 0 2
2 960 12 a001c 0 18 20030 558 959 1 0 2
2 961 12 a001c 0 18 20030 553 960 1 0 2
2 962 12 a001c 0 18 20030 548 961 1 0 2
2 963 12 a001c 0 18 20030 543 962 1 0 2
2 964 12 a001c 0 18 20030 538 963 1 0 2
2 965 12 a001c 0 18 20030 533 964 1 0 2
2 966 12 a001c 0 18 20030 528 965 1 0 2
2 967 12 a001c 0 18 20030 523 966 1 0 2
2 968 12 a001c 0 18 20030 518 967 1 0 2
2 969 12 a001c 0 18 20030 513 968 1 0 2
2 970 12 a001c 0 18 20030 508 969 1 0 2
2 971 12 a001c 0 18 20030 503 970 1 0 2
2 972 12 a001c 0 18 20030 498 971 1 0 2
2 973 12 a001c 0 18 20030 493 972 1 0 2
2 974 12 a001c 0 18 20030 488 973 1 0 2
2 975 12 a001c 0 18 20030 483 974 1 0 2
2 976 12 a001c 0 18 20030 478 975 1 0 2
2 977 12 a001c 0 18 20030 473 976 1 0 2
2 978 12 a001c 0 18 20030 468 977 1 0 2
2 979 11 d000d 0 1 10 0 0 c
2 980 11 90009 0 1 10 0 0 b
2 981 11 9000d 0 9 20030 979 980 1 0 2
2 982 11 8001d 0 8 20030 978 981 1 0 2
2 983 11 8001d 0 9 20030 463 982 1 0 2
2 984 11 30003 0 1 400 0 0 a
2 985 11 3001d 0 38 6022 983 984
2 986 9 110012 1 1 0 0 0 go
2 987 9 9000f 0 2a 20000 0 0 2 0 a
2 988 9 90012 2 27 21002 986 987 1 0 2
1 go 0 3 3000c 1 0 2
1 a 0 4 3000c 1 0 2
1 b 0 5 3000c 1 0 2
1 c 0 5 3000f 1 0 2
1 d 3 6 3000c 25 0 aa aa aa aa aa aa 2
1 e 0 7 3000c 1 0 2
4 985 988 988
4 988 985 0
*/

/* OUTPUT long_exp2.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : long_exp2.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp2.v                1/    1/    2       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           11:     a  <= ((( b  |  c ) & ...



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp2.v                0/   30/   30        0%             0/   30/   30        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 25'h000_0000
      ......................... 1->0: 25'h000_0000 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              long_exp2.v                         0/ 508/ 508        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    @(posedge  go)
                    |-----1------|

        Expression 1   (0/1)
        ^^^^^^^^^^^^^ - posedge
         * Event did not occur

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:     a  <= ((( b  |  c ) & 
                             |----1----|   
                            |------89-------
                           |------169-------
                    ((d[27:16] == 12'h0) && 
                     |--------2--------|    
                    |----------88------------
                    -----------89------------
                    -----------169-----------
                    (d[12:3] != 10'h0) && 
                    |-------3--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h1) && 
                    |-------4--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h2) && 
                    |-------5--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h3) && 
                    |-------6--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h4) && 
                    |-------7--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h5) && 
                    |-------8--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h6) && 
                    |-------9--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h7) && 
                    |-------10-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h8) && 
                    |-------11-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h9) && 
                    |-------12-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hA) && 
                    |-------13-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hB) && 
                    |-------14-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hC) && 
                    |-------15-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hD) && 
                    |-------16-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hE) && 
                    |-------17-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hF) && 
                    |-------18-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h10) && 
                    |-------19--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h11) && 
                    |-------20--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h12) && 
                    |-------21--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h13) && 
                    |-------22--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h14) && 
                    |-------23--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h15) && 
                    |-------24--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h16) && 
                    |-------25--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h17) && 
                    |-------26--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h18) && 
                    |-------27--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h19) && 
                    |-------28--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1A) && 
                    |-------29--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1B) && 
                    |-------30--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1C) && 
                    |-------31--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1D) && 
                    |-------32--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1E) && 
                    |-------33--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1F) && 
                    |-------34--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h20) && 
                    |-------35--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h21) && 
                    |-------36--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h22) && 
                    |-------37--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h23) && 
                    |-------38--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h24) && 
                    |-------39--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h25) && 
                    |-------40--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h26) && 
                    |-------41--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h27) && 
                    |-------42--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h28) && 
                    |-------43--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h29) && 
                    |-------44--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2A) && 
                    |-------45--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2B) && 
                    |-------46--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2C) && 
                    |-------47--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2D) && 
                    |-------48--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2E) && 
                    |-------49--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2F) && 
                    |-------50--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h30) && 
                    |-------51--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h31) && 
                    |-------52--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h32) && 
                    |-------53--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h33) && 
                    |-------54--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h34) && 
                    |-------55--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h35) && 
                    |-------56--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h36) && 
                    |-------57--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h37) && 
                    |-------58--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h38) && 
                    |-------59--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h39) && 
                    |-------60--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3A) && 
                    |-------61--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3B) && 
                    |-------62--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3C) && 
                    |-------63--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3D) && 
                    |-------64--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3E) && 
                    |-------65--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3F) && 
                    |-------66--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h40) && 
                    |-------67--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h41) && 
                    |-------68--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h42) && 
                    |-------69--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h43) && 
                    |-------70--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h44) && 
                    |-------71--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h45) && 
                    |-------72--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h46) && 
                    |-------73--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h47) && 
                    |-------74--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h48) && 
                    |-------75--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h49) && 
                    |-------76--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4A) && 
                    |-------77--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4B) && 
                    |-------78--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4C) && 
                    |-------79--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4D) && 
                    |-------80--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4E) && 
                    |-------81--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4F) && 
                    |-------82--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h50) && 
                    |-------83--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h51) && 
                    |-------84--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h52) && 
                    |-------85--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h53) && 
                    |-------86--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h54))) | 
                    |-------87--------|     
                    ---------88--------|    
                    ---------89---------|   
                    -----------169-----------
                    ( e  & 
                    |-168---
                    --169---
                    ((d[27:16] == 12'h0) && 
                     |-------90--------|    
                    |----------167-----------
                    -----------168-----------
                    -----------169-----------
                    (d[12:3] != 10'h0) && 
                    |-------91-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h1) && 
                    |-------92-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h2) && 
                    |-------93-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h3) && 
                    |-------94-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h4) && 
                    |-------95-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h5) && 
                    |-------96-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h6) && 
                    |-------97-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h7) && 
                    |-------98-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h8) && 
                    |-------99-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h9) && 
                    |------100-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hA) && 
                    |------101-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hB) && 
                    |------102-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hC) && 
                    |------103-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hD) && 
                    |------104-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hE) && 
                    |------105-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hF) && 
                    |------106-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h10) && 
                    |-------107-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h11) && 
                    |-------108-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h12) && 
                    |-------109-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h13) && 
                    |-------110-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h14) && 
                    |-------111-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h15) && 
                    |-------112-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h16) && 
                    |-------113-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h17) && 
                    |-------114-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h18) && 
                    |-------115-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h19) && 
                    |-------116-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1A) && 
                    |-------117-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1B) && 
                    |-------118-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1C) && 
                    |-------119-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1D) && 
                    |-------120-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1E) && 
                    |-------121-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1F) && 
                    |-------122-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h20) && 
                    |-------123-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h21) && 
                    |-------124-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h22) && 
                    |-------125-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h23) && 
                    |-------126-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h24) && 
                    |-------127-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h25) && 
                    |-------128-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h26) && 
                    |-------129-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h27) && 
                    |-------130-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h28) && 
                    |-------131-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h29) && 
                    |-------132-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2A) && 
                    |-------133-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2B) && 
                    |-------134-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2C) && 
                    |-------135-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2D) && 
                    |-------136-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2E) && 
                    |-------137-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2F) && 
                    |-------138-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h30) && 
                    |-------139-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h31) && 
                    |-------140-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h32) && 
                    |-------141-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h33) && 
                    |-------142-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h34) && 
                    |-------143-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h35) && 
                    |-------144-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h36) && 
                    |-------145-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h37) && 
                    |-------146-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h38) && 
                    |-------147-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h39) && 
                    |-------148-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3A) && 
                    |-------149-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3B) && 
                    |-------150-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3C) && 
                    |-------151-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3D) && 
                    |-------152-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3E) && 
                    |-------153-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3F) && 
                    |-------154-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h40) && 
                    |-------155-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h41) && 
                    |-------156-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h42) && 
                    |-------157-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h43) && 
                    |-------158-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h44) && 
                    |-------159-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h45) && 
                    |-------160-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h46) && 
                    |-------161-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h47) && 
                    |-------162-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h48) && 
                    |-------163-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h49) && 
                    |-------164-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h4A) && 
                    |-------165-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h4B))))
                    |-------166-------|   
                    --------167--------|  
                    ---------168--------| 
                    ---------169---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 3   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 4   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 5   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 6   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 7   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 8   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 9   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 10   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 11   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 12   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 13   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 14   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 15   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 16   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 17   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 18   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 19   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 20   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 21   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 22   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 23   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 24   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 25   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 26   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 27   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 28   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 29   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 30   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 31   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 32   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 33   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 34   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 35   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 36   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 37   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 38   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 39   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 40   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 41   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 42   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 43   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 44   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 45   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 46   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 47   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 48   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 49   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 50   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 51   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 52   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 53   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 54   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 55   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 56   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 57   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 58   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 59   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 60   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 61   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 62   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 63   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 64   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 65   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 66   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 67   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 68   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 69   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 70   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 71   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 72   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 73   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 74   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 75   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 76   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 77   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 78   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 79   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 80   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 81   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 82   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 83   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 84   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 85   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 86   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 87   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 88   (0/87)
        ^^^^^^^^^^^^^ - &&
         2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 | 16 | 17 | 18 | 19 | 20 | 21 | 22 | 23 | 24 |
        =0=|=0=|=0=|=0=|=0=|=0=|=0=|=0=|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *   *   *   *   *   *   *   *   *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         25 | 26 | 27 | 28 | 29 | 30 | 31 | 32 | 33 | 34 | 35 | 36 | 37 | 38 | 39 | 40 | 41 | 42 | 43 | 44 | 45 | 46 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         47 | 48 | 49 | 50 | 51 | 52 | 53 | 54 | 55 | 56 | 57 | 58 | 59 | 60 | 61 | 62 | 63 | 64 | 65 | 66 | 67 | 68 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         69 | 70 | 71 | 72 | 73 | 74 | 75 | 76 | 77 | 78 | 79 | 80 | 81 | 82 | 83 | 84 | 85 | 86 | 87 | All
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|==1==
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *     *  

        Expression 89   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 90   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 91   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 92   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 93   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 94   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 95   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 96   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 97   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 98   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 99   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 100   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 101   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 102   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 103   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 104   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 105   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 106   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 107   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 108   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 109   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 110   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 111   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 112   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 113   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 114   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 115   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 116   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 117   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 118   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 119   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 120   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 121   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 122   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 123   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 124   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 125   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 126   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 127   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 128   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 129   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 130   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 131   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 132   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 133   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 134   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 135   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 136   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 137   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 138   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 139   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 140   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 141   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 142   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 143   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 144   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 145   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 146   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 147   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 148   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 149   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 150   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 151   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 152   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 153   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 154   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 155   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 156   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 157   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 158   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 159   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 160   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 161   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 162   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 163   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 164   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 165   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 166   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 167   (0/78)
        ^^^^^^^^^^^^^ - &&
         90 | 91 | 92 | 93 | 94 | 95 | 96 | 97 | 98 | 99 | 100 | 101 | 102 | 103 | 104 | 105 | 106 | 107 | 108 | 109 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *    *    *    *    *    *    *    *    *    *    *     *     *     *     *     *     *     *     *     *    

         110 | 111 | 112 | 113 | 114 | 115 | 116 | 117 | 118 | 119 | 120 | 121 | 122 | 123 | 124 | 125 | 126 | 127 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         128 | 129 | 130 | 131 | 132 | 133 | 134 | 135 | 136 | 137 | 138 | 139 | 140 | 141 | 142 | 143 | 144 | 145 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         146 | 147 | 148 | 149 | 150 | 151 | 152 | 153 | 154 | 155 | 156 | 157 | 158 | 159 | 160 | 161 | 162 | 163 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         164 | 165 | 166 | All
        =0===|=0===|=0===|==1==
         *     *     *      *  

        Expression 168   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 169   (0/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp2.v               0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT long_exp2.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : long_exp2.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp2.v                1/    1/    2       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           11:     a  <= ((( b  |  c ) & ...



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp2.v                0/   30/   30        0%             0/   30/   30        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 25'h000_0000
      ......................... 1->0: 25'h000_0000 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              long_exp2.v                         0/ 508/ 508        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    @(posedge  go)
                    |-----1------|

        Expression 1   (0/1)
        ^^^^^^^^^^^^^ - posedge
         * Event did not occur

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:     a  <= ((( b  |  c ) & 
                             |----1----|   
                            |------89-------
                           |------169-------
                    ((d[27:16] == 12'h0) && (d[12:3] != 10'h0) && (d[12:3] != 10'h1) && (d[12:3] != 10'h2) && 
                     |--------2--------|    |-------3--------|    |-------4--------|    |-------5--------|    
                    |-------------------------------------------88---------------------------------------------
                    --------------------------------------------89---------------------------------------------
                    --------------------------------------------169--------------------------------------------
                    (d[12:3] != 10'h3) && (d[12:3] != 10'h4) && (d[12:3] != 10'h5) && (d[12:3] != 10'h6) && 
                    |-------6--------|    |-------7--------|    |-------8--------|    |-------9--------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'h7) && (d[12:3] != 10'h8) && (d[12:3] != 10'h9) && (d[12:3] != 10'hA) && 
                    |-------10-------|    |-------11-------|    |-------12-------|    |-------13-------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hB) && (d[12:3] != 10'hC) && (d[12:3] != 10'hD) && (d[12:3] != 10'hE) && 
                    |-------14-------|    |-------15-------|    |-------16-------|    |-------17-------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hF) && (d[12:3] != 10'h10) && (d[12:3] != 10'h11) && (d[12:3] != 10'h12) && 
                    |-------18-------|    |-------19--------|    |-------20--------|    |-------21--------|    
                    ---------------------------------------------88---------------------------------------------
                    ---------------------------------------------89---------------------------------------------
                    --------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h13) && (d[12:3] != 10'h14) && (d[12:3] != 10'h15) && (d[12:3] != 10'h16) && 
                    |-------22--------|    |-------23--------|    |-------24--------|    |-------25--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h17) && (d[12:3] != 10'h18) && (d[12:3] != 10'h19) && (d[12:3] != 10'h1A) && 
                    |-------26--------|    |-------27--------|    |-------28--------|    |-------29--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1B) && (d[12:3] != 10'h1C) && (d[12:3] != 10'h1D) && (d[12:3] != 10'h1E) && 
                    |-------30--------|    |-------31--------|    |-------32--------|    |-------33--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1F) && (d[12:3] != 10'h20) && (d[12:3] != 10'h21) && (d[12:3] != 10'h22) && 
                    |-------34--------|    |-------35--------|    |-------36--------|    |-------37--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h23) && (d[12:3] != 10'h24) && (d[12:3] != 10'h25) && (d[12:3] != 10'h26) && 
                    |-------38--------|    |-------39--------|    |-------40--------|    |-------41--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h27) && (d[12:3] != 10'h28) && (d[12:3] != 10'h29) && (d[12:3] != 10'h2A) && 
                    |-------42--------|    |-------43--------|    |-------44--------|    |-------45--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2B) && (d[12:3] != 10'h2C) && (d[12:3] != 10'h2D) && (d[12:3] != 10'h2E) && 
                    |-------46--------|    |-------47--------|    |-------48--------|    |-------49--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2F) && (d[12:3] != 10'h30) && (d[12:3] != 10'h31) && (d[12:3] != 10'h32) && 
                    |-------50--------|    |-------51--------|    |-------52--------|    |-------53--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h33) && (d[12:3] != 10'h34) && (d[12:3] != 10'h35) && (d[12:3] != 10'h36) && 
                    |-------54--------|    |-------55--------|    |-------56--------|    |-------57--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h37) && (d[12:3] != 10'h38) && (d[12:3] != 10'h39) && (d[12:3] != 10'h3A) && 
                    |-------58--------|    |-------59--------|    |-------60--------|    |-------61--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3B) && (d[12:3] != 10'h3C) && (d[12:3] != 10'h3D) && (d[12:3] != 10'h3E) && 
                    |-------62--------|    |-------63--------|    |-------64--------|    |-------65--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3F) && (d[12:3] != 10'h40) && (d[12:3] != 10'h41) && (d[12:3] != 10'h42) && 
                    |-------66--------|    |-------67--------|    |-------68--------|    |-------69--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h43) && (d[12:3] != 10'h44) && (d[12:3] != 10'h45) && (d[12:3] != 10'h46) && 
                    |-------70--------|    |-------71--------|    |-------72--------|    |-------73--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h47) && (d[12:3] != 10'h48) && (d[12:3] != 10'h49) && (d[12:3] != 10'h4A) && 
                    |-------74--------|    |-------75--------|    |-------76--------|    |-------77--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4B) && (d[12:3] != 10'h4C) && (d[12:3] != 10'h4D) && (d[12:3] != 10'h4E) && 
                    |-------78--------|    |-------79--------|    |-------80--------|    |-------81--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4F) && (d[12:3] != 10'h50) && (d[12:3] != 10'h51) && (d[12:3] != 10'h52) && 
                    |-------82--------|    |-------83--------|    |-------84--------|    |-------85--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h53) && (d[12:3] != 10'h54))) | 
                    |-------86--------|    |-------87--------|     
                    --------------------88--------------------|    
                    ---------------------89--------------------|   
                    ----------------------169-----------------------
                    ( e  & ((d[27:16] == 12'h0) && (d[12:3] != 10'h0) && (d[12:3] != 10'h1) && (d[12:3] != 10'h2) && 
                            |-------90--------|    |-------91-------|    |-------92-------|    |-------93-------|    
                           |-------------------------------------------167--------------------------------------------
                    |----------------------------------------------168------------------------------------------------
                    -----------------------------------------------169------------------------------------------------
                    (d[12:3] != 10'h3) && (d[12:3] != 10'h4) && (d[12:3] != 10'h5) && (d[12:3] != 10'h6) && 
                    |-------94-------|    |-------95-------|    |-------96-------|    |-------97-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'h7) && (d[12:3] != 10'h8) && (d[12:3] != 10'h9) && (d[12:3] != 10'hA) && 
                    |-------98-------|    |-------99-------|    |------100-------|    |------101-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hB) && (d[12:3] != 10'hC) && (d[12:3] != 10'hD) && (d[12:3] != 10'hE) && 
                    |------102-------|    |------103-------|    |------104-------|    |------105-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hF) && (d[12:3] != 10'h10) && (d[12:3] != 10'h11) && (d[12:3] != 10'h12) && 
                    |------106-------|    |-------107-------|    |-------108-------|    |-------109-------|    
                    --------------------------------------------167---------------------------------------------
                    --------------------------------------------168---------------------------------------------
                    --------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h13) && (d[12:3] != 10'h14) && (d[12:3] != 10'h15) && (d[12:3] != 10'h16) && 
                    |-------110-------|    |-------111-------|    |-------112-------|    |-------113-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h17) && (d[12:3] != 10'h18) && (d[12:3] != 10'h19) && (d[12:3] != 10'h1A) && 
                    |-------114-------|    |-------115-------|    |-------116-------|    |-------117-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1B) && (d[12:3] != 10'h1C) && (d[12:3] != 10'h1D) && (d[12:3] != 10'h1E) && 
                    |-------118-------|    |-------119-------|    |-------120-------|    |-------121-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1F) && (d[12:3] != 10'h20) && (d[12:3] != 10'h21) && (d[12:3] != 10'h22) && 
                    |-------122-------|    |-------123-------|    |-------124-------|    |-------125-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h23) && (d[12:3] != 10'h24) && (d[12:3] != 10'h25) && (d[12:3] != 10'h26) && 
                    |-------126-------|    |-------127-------|    |-------128-------|    |-------129-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h27) && (d[12:3] != 10'h28) && (d[12:3] != 10'h29) && (d[12:3] != 10'h2A) && 
                    |-------130-------|    |-------131-------|    |-------132-------|    |-------133-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2B) && (d[12:3] != 10'h2C) && (d[12:3] != 10'h2D) && (d[12:3] != 10'h2E) && 
                    |-------134-------|    |-------135-------|    |-------136-------|    |-------137-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2F) && (d[12:3] != 10'h30) && (d[12:3] != 10'h31) && (d[12:3] != 10'h32) && 
                    |-------138-------|    |-------139-------|    |-------140-------|    |-------141-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h33) && (d[12:3] != 10'h34) && (d[12:3] != 10'h35) && (d[12:3] != 10'h36) && 
                    |-------142-------|    |-------143-------|    |-------144-------|    |-------145-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h37) && (d[12:3] != 10'h38) && (d[12:3] != 10'h39) && (d[12:3] != 10'h3A) && 
                    |-------146-------|    |-------147-------|    |-------148-------|    |-------149-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3B) && (d[12:3] != 10'h3C) && (d[12:3] != 10'h3D) && (d[12:3] != 10'h3E) && 
                    |-------150-------|    |-------151-------|    |-------152-------|    |-------153-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3F) && (d[12:3] != 10'h40) && (d[12:3] != 10'h41) && (d[12:3] != 10'h42) && 
                    |-------154-------|    |-------155-------|    |-------156-------|    |-------157-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h43) && (d[12:3] != 10'h44) && (d[12:3] != 10'h45) && (d[12:3] != 10'h46) && 
                    |-------158-------|    |-------159-------|    |-------160-------|    |-------161-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h47) && (d[12:3] != 10'h48) && (d[12:3] != 10'h49) && (d[12:3] != 10'h4A) && 
                    |-------162-------|    |-------163-------|    |-------164-------|    |-------165-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4B))))
                    |-------166-------|   
                    --------167--------|  
                    ---------168--------| 
                    ---------169---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 3   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 4   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 5   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 6   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 7   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 8   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 9   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 10   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 11   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 12   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 13   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 14   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 15   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 16   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 17   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 18   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 19   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 20   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 21   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 22   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 23   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 24   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 25   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 26   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 27   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 28   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 29   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 30   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 31   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 32   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 33   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 34   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 35   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 36   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 37   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 38   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 39   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 40   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 41   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 42   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 43   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 44   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 45   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 46   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 47   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 48   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 49   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 50   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 51   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 52   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 53   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 54   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 55   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 56   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 57   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 58   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 59   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 60   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 61   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 62   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 63   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 64   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 65   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 66   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 67   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 68   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 69   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 70   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 71   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 72   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 73   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 74   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 75   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 76   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 77   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 78   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 79   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 80   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 81   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 82   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 83   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 84   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 85   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 86   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 87   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 88   (0/87)
        ^^^^^^^^^^^^^ - &&
         2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 | 16 | 17 | 18 | 19 | 20 | 21 | 22 | 23 | 24 |
        =0=|=0=|=0=|=0=|=0=|=0=|=0=|=0=|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *   *   *   *   *   *   *   *   *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         25 | 26 | 27 | 28 | 29 | 30 | 31 | 32 | 33 | 34 | 35 | 36 | 37 | 38 | 39 | 40 | 41 | 42 | 43 | 44 | 45 | 46 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         47 | 48 | 49 | 50 | 51 | 52 | 53 | 54 | 55 | 56 | 57 | 58 | 59 | 60 | 61 | 62 | 63 | 64 | 65 | 66 | 67 | 68 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         69 | 70 | 71 | 72 | 73 | 74 | 75 | 76 | 77 | 78 | 79 | 80 | 81 | 82 | 83 | 84 | 85 | 86 | 87 | All
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|==1==
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *     *  

        Expression 89   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 90   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 91   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 92   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 93   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 94   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 95   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 96   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 97   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 98   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 99   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 100   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 101   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 102   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 103   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 104   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 105   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 106   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 107   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 108   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 109   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 110   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 111   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 112   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 113   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 114   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 115   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 116   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 117   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 118   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 119   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 120   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 121   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 122   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 123   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 124   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 125   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 126   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 127   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 128   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 129   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 130   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 131   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 132   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 133   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 134   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 135   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 136   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 137   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 138   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 139   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 140   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 141   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 142   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 143   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 144   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 145   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 146   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 147   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 148   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 149   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 150   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 151   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 152   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 153   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 154   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 155   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 156   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 157   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 158   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 159   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 160   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 161   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 162   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 163   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 164   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 165   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 166   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 167   (0/78)
        ^^^^^^^^^^^^^ - &&
         90 | 91 | 92 | 93 | 94 | 95 | 96 | 97 | 98 | 99 | 100 | 101 | 102 | 103 | 104 | 105 | 106 | 107 | 108 | 109 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *    *    *    *    *    *    *    *    *    *    *     *     *     *     *     *     *     *     *     *    

         110 | 111 | 112 | 113 | 114 | 115 | 116 | 117 | 118 | 119 | 120 | 121 | 122 | 123 | 124 | 125 | 126 | 127 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         128 | 129 | 130 | 131 | 132 | 133 | 134 | 135 | 136 | 137 | 138 | 139 | 140 | 141 | 142 | 143 | 144 | 145 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         146 | 147 | 148 | 149 | 150 | 151 | 152 | 153 | 154 | 155 | 156 | 157 | 158 | 159 | 160 | 161 | 162 | 163 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         164 | 165 | 166 | All
        =0===|=0===|=0===|==1==
         *     *     *      *  

        Expression 168   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 169   (0/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    long_exp2.v               0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT long_exp2.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : long_exp2.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/    1/    2       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           11:     a  <= ((( b  |  c ) & ...



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/   30/   30        0%             0/   30/   30        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 25'h000_0000
      ......................... 1->0: 25'h000_0000 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/ 508/ 508        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    @(posedge  go)
                    |-----1------|

        Expression 1   (0/1)
        ^^^^^^^^^^^^^ - posedge
         * Event did not occur

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:     a  <= ((( b  |  c ) & 
                             |----1----|   
                            |------89-------
                           |------169-------
                    ((d[27:16] == 12'h0) && 
                     |--------2--------|    
                    |----------88------------
                    -----------89------------
                    -----------169-----------
                    (d[12:3] != 10'h0) && 
                    |-------3--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h1) && 
                    |-------4--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h2) && 
                    |-------5--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h3) && 
                    |-------6--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h4) && 
                    |-------7--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h5) && 
                    |-------8--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h6) && 
                    |-------9--------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h7) && 
                    |-------10-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h8) && 
                    |-------11-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h9) && 
                    |-------12-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hA) && 
                    |-------13-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hB) && 
                    |-------14-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hC) && 
                    |-------15-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hD) && 
                    |-------16-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hE) && 
                    |-------17-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'hF) && 
                    |-------18-------|    
                    ----------88-----------
                    ----------89-----------
                    ----------169----------
                    (d[12:3] != 10'h10) && 
                    |-------19--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h11) && 
                    |-------20--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h12) && 
                    |-------21--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h13) && 
                    |-------22--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h14) && 
                    |-------23--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h15) && 
                    |-------24--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h16) && 
                    |-------25--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h17) && 
                    |-------26--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h18) && 
                    |-------27--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h19) && 
                    |-------28--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1A) && 
                    |-------29--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1B) && 
                    |-------30--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1C) && 
                    |-------31--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1D) && 
                    |-------32--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1E) && 
                    |-------33--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h1F) && 
                    |-------34--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h20) && 
                    |-------35--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h21) && 
                    |-------36--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h22) && 
                    |-------37--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h23) && 
                    |-------38--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h24) && 
                    |-------39--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h25) && 
                    |-------40--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h26) && 
                    |-------41--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h27) && 
                    |-------42--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h28) && 
                    |-------43--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h29) && 
                    |-------44--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2A) && 
                    |-------45--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2B) && 
                    |-------46--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2C) && 
                    |-------47--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2D) && 
                    |-------48--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2E) && 
                    |-------49--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h2F) && 
                    |-------50--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h30) && 
                    |-------51--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h31) && 
                    |-------52--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h32) && 
                    |-------53--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h33) && 
                    |-------54--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h34) && 
                    |-------55--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h35) && 
                    |-------56--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h36) && 
                    |-------57--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h37) && 
                    |-------58--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h38) && 
                    |-------59--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h39) && 
                    |-------60--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3A) && 
                    |-------61--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3B) && 
                    |-------62--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3C) && 
                    |-------63--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3D) && 
                    |-------64--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3E) && 
                    |-------65--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h3F) && 
                    |-------66--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h40) && 
                    |-------67--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h41) && 
                    |-------68--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h42) && 
                    |-------69--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h43) && 
                    |-------70--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h44) && 
                    |-------71--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h45) && 
                    |-------72--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h46) && 
                    |-------73--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h47) && 
                    |-------74--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h48) && 
                    |-------75--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h49) && 
                    |-------76--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4A) && 
                    |-------77--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4B) && 
                    |-------78--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4C) && 
                    |-------79--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4D) && 
                    |-------80--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4E) && 
                    |-------81--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h4F) && 
                    |-------82--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h50) && 
                    |-------83--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h51) && 
                    |-------84--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h52) && 
                    |-------85--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h53) && 
                    |-------86--------|    
                    -----------88-----------
                    -----------89-----------
                    ----------169-----------
                    (d[12:3] != 10'h54))) | 
                    |-------87--------|     
                    ---------88--------|    
                    ---------89---------|   
                    -----------169-----------
                    ( e  & 
                    |-168---
                    --169---
                    ((d[27:16] == 12'h0) && 
                     |-------90--------|    
                    |----------167-----------
                    -----------168-----------
                    -----------169-----------
                    (d[12:3] != 10'h0) && 
                    |-------91-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h1) && 
                    |-------92-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h2) && 
                    |-------93-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h3) && 
                    |-------94-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h4) && 
                    |-------95-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h5) && 
                    |-------96-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h6) && 
                    |-------97-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h7) && 
                    |-------98-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h8) && 
                    |-------99-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h9) && 
                    |------100-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hA) && 
                    |------101-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hB) && 
                    |------102-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hC) && 
                    |------103-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hD) && 
                    |------104-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hE) && 
                    |------105-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'hF) && 
                    |------106-------|    
                    ----------167----------
                    ----------168----------
                    ----------169----------
                    (d[12:3] != 10'h10) && 
                    |-------107-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h11) && 
                    |-------108-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h12) && 
                    |-------109-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h13) && 
                    |-------110-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h14) && 
                    |-------111-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h15) && 
                    |-------112-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h16) && 
                    |-------113-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h17) && 
                    |-------114-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h18) && 
                    |-------115-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h19) && 
                    |-------116-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1A) && 
                    |-------117-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1B) && 
                    |-------118-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1C) && 
                    |-------119-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1D) && 
                    |-------120-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1E) && 
                    |-------121-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h1F) && 
                    |-------122-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h20) && 
                    |-------123-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h21) && 
                    |-------124-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h22) && 
                    |-------125-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h23) && 
                    |-------126-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h24) && 
                    |-------127-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h25) && 
                    |-------128-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h26) && 
                    |-------129-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h27) && 
                    |-------130-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h28) && 
                    |-------131-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h29) && 
                    |-------132-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2A) && 
                    |-------133-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2B) && 
                    |-------134-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2C) && 
                    |-------135-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2D) && 
                    |-------136-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2E) && 
                    |-------137-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h2F) && 
                    |-------138-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h30) && 
                    |-------139-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h31) && 
                    |-------140-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h32) && 
                    |-------141-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h33) && 
                    |-------142-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h34) && 
                    |-------143-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h35) && 
                    |-------144-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h36) && 
                    |-------145-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h37) && 
                    |-------146-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h38) && 
                    |-------147-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h39) && 
                    |-------148-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3A) && 
                    |-------149-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3B) && 
                    |-------150-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3C) && 
                    |-------151-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3D) && 
                    |-------152-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3E) && 
                    |-------153-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h3F) && 
                    |-------154-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h40) && 
                    |-------155-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h41) && 
                    |-------156-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h42) && 
                    |-------157-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h43) && 
                    |-------158-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h44) && 
                    |-------159-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h45) && 
                    |-------160-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h46) && 
                    |-------161-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h47) && 
                    |-------162-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h48) && 
                    |-------163-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h49) && 
                    |-------164-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h4A) && 
                    |-------165-------|    
                    ----------167-----------
                    ----------168-----------
                    ----------169-----------
                    (d[12:3] != 10'h4B))))
                    |-------166-------|   
                    --------167--------|  
                    ---------168--------| 
                    ---------169---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 3   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 4   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 5   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 6   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 7   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 8   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 9   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 10   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 11   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 12   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 13   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 14   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 15   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 16   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 17   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 18   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 19   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 20   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 21   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 22   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 23   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 24   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 25   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 26   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 27   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 28   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 29   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 30   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 31   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 32   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 33   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 34   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 35   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 36   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 37   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 38   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 39   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 40   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 41   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 42   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 43   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 44   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 45   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 46   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 47   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 48   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 49   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 50   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 51   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 52   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 53   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 54   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 55   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 56   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 57   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 58   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 59   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 60   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 61   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 62   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 63   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 64   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 65   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 66   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 67   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 68   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 69   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 70   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 71   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 72   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 73   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 74   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 75   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 76   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 77   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 78   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 79   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 80   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 81   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 82   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 83   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 84   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 85   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 86   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 87   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 88   (0/87)
        ^^^^^^^^^^^^^ - &&
         2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 | 16 | 17 | 18 | 19 | 20 | 21 | 22 | 23 | 24 |
        =0=|=0=|=0=|=0=|=0=|=0=|=0=|=0=|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *   *   *   *   *   *   *   *   *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         25 | 26 | 27 | 28 | 29 | 30 | 31 | 32 | 33 | 34 | 35 | 36 | 37 | 38 | 39 | 40 | 41 | 42 | 43 | 44 | 45 | 46 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         47 | 48 | 49 | 50 | 51 | 52 | 53 | 54 | 55 | 56 | 57 | 58 | 59 | 60 | 61 | 62 | 63 | 64 | 65 | 66 | 67 | 68 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         69 | 70 | 71 | 72 | 73 | 74 | 75 | 76 | 77 | 78 | 79 | 80 | 81 | 82 | 83 | 84 | 85 | 86 | 87 | All
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|==1==
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *     *  

        Expression 89   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 90   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 91   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 92   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 93   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 94   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 95   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 96   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 97   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 98   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 99   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 100   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 101   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 102   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 103   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 104   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 105   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 106   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 107   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 108   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 109   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 110   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 111   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 112   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 113   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 114   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 115   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 116   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 117   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 118   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 119   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 120   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 121   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 122   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 123   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 124   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 125   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 126   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 127   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 128   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 129   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 130   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 131   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 132   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 133   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 134   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 135   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 136   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 137   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 138   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 139   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 140   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 141   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 142   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 143   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 144   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 145   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 146   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 147   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 148   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 149   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 150   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 151   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 152   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 153   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 154   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 155   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 156   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 157   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 158   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 159   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 160   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 161   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 162   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 163   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 164   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 165   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 166   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 167   (0/78)
        ^^^^^^^^^^^^^ - &&
         90 | 91 | 92 | 93 | 94 | 95 | 96 | 97 | 98 | 99 | 100 | 101 | 102 | 103 | 104 | 105 | 106 | 107 | 108 | 109 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *    *    *    *    *    *    *    *    *    *    *     *     *     *     *     *     *     *     *     *    

         110 | 111 | 112 | 113 | 114 | 115 | 116 | 117 | 118 | 119 | 120 | 121 | 122 | 123 | 124 | 125 | 126 | 127 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         128 | 129 | 130 | 131 | 132 | 133 | 134 | 135 | 136 | 137 | 138 | 139 | 140 | 141 | 142 | 143 | 144 | 145 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         146 | 147 | 148 | 149 | 150 | 151 | 152 | 153 | 154 | 155 | 156 | 157 | 158 | 159 | 160 | 161 | 162 | 163 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         164 | 165 | 166 | All
        =0===|=0===|=0===|==1==
         *     *     *      *  

        Expression 168   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 169   (0/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT long_exp2.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : long_exp2.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/    1/    2       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           11:     a  <= ((( b  |  c ) & ...



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/   30/   30        0%             0/   30/   30        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      go                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 25'h000_0000
      ......................... 1->0: 25'h000_0000 ...
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/ 508/ 508        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: long_exp2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    @(posedge  go)
                    |-----1------|

        Expression 1   (0/1)
        ^^^^^^^^^^^^^ - posedge
         * Event did not occur

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:     a  <= ((( b  |  c ) & 
                             |----1----|   
                            |------89-------
                           |------169-------
                    ((d[27:16] == 12'h0) && (d[12:3] != 10'h0) && (d[12:3] != 10'h1) && (d[12:3] != 10'h2) && 
                     |--------2--------|    |-------3--------|    |-------4--------|    |-------5--------|    
                    |-------------------------------------------88---------------------------------------------
                    --------------------------------------------89---------------------------------------------
                    --------------------------------------------169--------------------------------------------
                    (d[12:3] != 10'h3) && (d[12:3] != 10'h4) && (d[12:3] != 10'h5) && (d[12:3] != 10'h6) && 
                    |-------6--------|    |-------7--------|    |-------8--------|    |-------9--------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'h7) && (d[12:3] != 10'h8) && (d[12:3] != 10'h9) && (d[12:3] != 10'hA) && 
                    |-------10-------|    |-------11-------|    |-------12-------|    |-------13-------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hB) && (d[12:3] != 10'hC) && (d[12:3] != 10'hD) && (d[12:3] != 10'hE) && 
                    |-------14-------|    |-------15-------|    |-------16-------|    |-------17-------|    
                    -------------------------------------------88--------------------------------------------
                    -------------------------------------------89--------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hF) && (d[12:3] != 10'h10) && (d[12:3] != 10'h11) && (d[12:3] != 10'h12) && 
                    |-------18-------|    |-------19--------|    |-------20--------|    |-------21--------|    
                    ---------------------------------------------88---------------------------------------------
                    ---------------------------------------------89---------------------------------------------
                    --------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h13) && (d[12:3] != 10'h14) && (d[12:3] != 10'h15) && (d[12:3] != 10'h16) && 
                    |-------22--------|    |-------23--------|    |-------24--------|    |-------25--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h17) && (d[12:3] != 10'h18) && (d[12:3] != 10'h19) && (d[12:3] != 10'h1A) && 
                    |-------26--------|    |-------27--------|    |-------28--------|    |-------29--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1B) && (d[12:3] != 10'h1C) && (d[12:3] != 10'h1D) && (d[12:3] != 10'h1E) && 
                    |-------30--------|    |-------31--------|    |-------32--------|    |-------33--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1F) && (d[12:3] != 10'h20) && (d[12:3] != 10'h21) && (d[12:3] != 10'h22) && 
                    |-------34--------|    |-------35--------|    |-------36--------|    |-------37--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h23) && (d[12:3] != 10'h24) && (d[12:3] != 10'h25) && (d[12:3] != 10'h26) && 
                    |-------38--------|    |-------39--------|    |-------40--------|    |-------41--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h27) && (d[12:3] != 10'h28) && (d[12:3] != 10'h29) && (d[12:3] != 10'h2A) && 
                    |-------42--------|    |-------43--------|    |-------44--------|    |-------45--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2B) && (d[12:3] != 10'h2C) && (d[12:3] != 10'h2D) && (d[12:3] != 10'h2E) && 
                    |-------46--------|    |-------47--------|    |-------48--------|    |-------49--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2F) && (d[12:3] != 10'h30) && (d[12:3] != 10'h31) && (d[12:3] != 10'h32) && 
                    |-------50--------|    |-------51--------|    |-------52--------|    |-------53--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h33) && (d[12:3] != 10'h34) && (d[12:3] != 10'h35) && (d[12:3] != 10'h36) && 
                    |-------54--------|    |-------55--------|    |-------56--------|    |-------57--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h37) && (d[12:3] != 10'h38) && (d[12:3] != 10'h39) && (d[12:3] != 10'h3A) && 
                    |-------58--------|    |-------59--------|    |-------60--------|    |-------61--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3B) && (d[12:3] != 10'h3C) && (d[12:3] != 10'h3D) && (d[12:3] != 10'h3E) && 
                    |-------62--------|    |-------63--------|    |-------64--------|    |-------65--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3F) && (d[12:3] != 10'h40) && (d[12:3] != 10'h41) && (d[12:3] != 10'h42) && 
                    |-------66--------|    |-------67--------|    |-------68--------|    |-------69--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h43) && (d[12:3] != 10'h44) && (d[12:3] != 10'h45) && (d[12:3] != 10'h46) && 
                    |-------70--------|    |-------71--------|    |-------72--------|    |-------73--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h47) && (d[12:3] != 10'h48) && (d[12:3] != 10'h49) && (d[12:3] != 10'h4A) && 
                    |-------74--------|    |-------75--------|    |-------76--------|    |-------77--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4B) && (d[12:3] != 10'h4C) && (d[12:3] != 10'h4D) && (d[12:3] != 10'h4E) && 
                    |-------78--------|    |-------79--------|    |-------80--------|    |-------81--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4F) && (d[12:3] != 10'h50) && (d[12:3] != 10'h51) && (d[12:3] != 10'h52) && 
                    |-------82--------|    |-------83--------|    |-------84--------|    |-------85--------|    
                    ---------------------------------------------88----------------------------------------------
                    ---------------------------------------------89----------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h53) && (d[12:3] != 10'h54))) | 
                    |-------86--------|    |-------87--------|     
                    --------------------88--------------------|    
                    ---------------------89--------------------|   
                    ----------------------169-----------------------
                    ( e  & ((d[27:16] == 12'h0) && (d[12:3] != 10'h0) && (d[12:3] != 10'h1) && (d[12:3] != 10'h2) && 
                            |-------90--------|    |-------91-------|    |-------92-------|    |-------93-------|    
                           |-------------------------------------------167--------------------------------------------
                    |----------------------------------------------168------------------------------------------------
                    -----------------------------------------------169------------------------------------------------
                    (d[12:3] != 10'h3) && (d[12:3] != 10'h4) && (d[12:3] != 10'h5) && (d[12:3] != 10'h6) && 
                    |-------94-------|    |-------95-------|    |-------96-------|    |-------97-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'h7) && (d[12:3] != 10'h8) && (d[12:3] != 10'h9) && (d[12:3] != 10'hA) && 
                    |-------98-------|    |-------99-------|    |------100-------|    |------101-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hB) && (d[12:3] != 10'hC) && (d[12:3] != 10'hD) && (d[12:3] != 10'hE) && 
                    |------102-------|    |------103-------|    |------104-------|    |------105-------|    
                    -------------------------------------------167-------------------------------------------
                    -------------------------------------------168-------------------------------------------
                    -------------------------------------------169-------------------------------------------
                    (d[12:3] != 10'hF) && (d[12:3] != 10'h10) && (d[12:3] != 10'h11) && (d[12:3] != 10'h12) && 
                    |------106-------|    |-------107-------|    |-------108-------|    |-------109-------|    
                    --------------------------------------------167---------------------------------------------
                    --------------------------------------------168---------------------------------------------
                    --------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h13) && (d[12:3] != 10'h14) && (d[12:3] != 10'h15) && (d[12:3] != 10'h16) && 
                    |-------110-------|    |-------111-------|    |-------112-------|    |-------113-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h17) && (d[12:3] != 10'h18) && (d[12:3] != 10'h19) && (d[12:3] != 10'h1A) && 
                    |-------114-------|    |-------115-------|    |-------116-------|    |-------117-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1B) && (d[12:3] != 10'h1C) && (d[12:3] != 10'h1D) && (d[12:3] != 10'h1E) && 
                    |-------118-------|    |-------119-------|    |-------120-------|    |-------121-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h1F) && (d[12:3] != 10'h20) && (d[12:3] != 10'h21) && (d[12:3] != 10'h22) && 
                    |-------122-------|    |-------123-------|    |-------124-------|    |-------125-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h23) && (d[12:3] != 10'h24) && (d[12:3] != 10'h25) && (d[12:3] != 10'h26) && 
                    |-------126-------|    |-------127-------|    |-------128-------|    |-------129-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h27) && (d[12:3] != 10'h28) && (d[12:3] != 10'h29) && (d[12:3] != 10'h2A) && 
                    |-------130-------|    |-------131-------|    |-------132-------|    |-------133-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2B) && (d[12:3] != 10'h2C) && (d[12:3] != 10'h2D) && (d[12:3] != 10'h2E) && 
                    |-------134-------|    |-------135-------|    |-------136-------|    |-------137-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h2F) && (d[12:3] != 10'h30) && (d[12:3] != 10'h31) && (d[12:3] != 10'h32) && 
                    |-------138-------|    |-------139-------|    |-------140-------|    |-------141-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h33) && (d[12:3] != 10'h34) && (d[12:3] != 10'h35) && (d[12:3] != 10'h36) && 
                    |-------142-------|    |-------143-------|    |-------144-------|    |-------145-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h37) && (d[12:3] != 10'h38) && (d[12:3] != 10'h39) && (d[12:3] != 10'h3A) && 
                    |-------146-------|    |-------147-------|    |-------148-------|    |-------149-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3B) && (d[12:3] != 10'h3C) && (d[12:3] != 10'h3D) && (d[12:3] != 10'h3E) && 
                    |-------150-------|    |-------151-------|    |-------152-------|    |-------153-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h3F) && (d[12:3] != 10'h40) && (d[12:3] != 10'h41) && (d[12:3] != 10'h42) && 
                    |-------154-------|    |-------155-------|    |-------156-------|    |-------157-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h43) && (d[12:3] != 10'h44) && (d[12:3] != 10'h45) && (d[12:3] != 10'h46) && 
                    |-------158-------|    |-------159-------|    |-------160-------|    |-------161-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h47) && (d[12:3] != 10'h48) && (d[12:3] != 10'h49) && (d[12:3] != 10'h4A) && 
                    |-------162-------|    |-------163-------|    |-------164-------|    |-------165-------|    
                    ---------------------------------------------167---------------------------------------------
                    ---------------------------------------------168---------------------------------------------
                    ---------------------------------------------169---------------------------------------------
                    (d[12:3] != 10'h4B))))
                    |-------166-------|   
                    --------167--------|  
                    ---------168--------| 
                    ---------169---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 3   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 4   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 5   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 6   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 7   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 8   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 9   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 10   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 11   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 12   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 13   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 14   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 15   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 16   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 17   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 18   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 19   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 20   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 21   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 22   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 23   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 24   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 25   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 26   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 27   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 28   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 29   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 30   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 31   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 32   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 33   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 34   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 35   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 36   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 37   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 38   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 39   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 40   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 41   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 42   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 43   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 44   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 45   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 46   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 47   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 48   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 49   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 50   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 51   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 52   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 53   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 54   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 55   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 56   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 57   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 58   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 59   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 60   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 61   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 62   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 63   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 64   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 65   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 66   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 67   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 68   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 69   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 70   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 71   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 72   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 73   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 74   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 75   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 76   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 77   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 78   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 79   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 80   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 81   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 82   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 83   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 84   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 85   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 86   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 87   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 88   (0/87)
        ^^^^^^^^^^^^^ - &&
         2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 | 16 | 17 | 18 | 19 | 20 | 21 | 22 | 23 | 24 |
        =0=|=0=|=0=|=0=|=0=|=0=|=0=|=0=|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *   *   *   *   *   *   *   *   *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         25 | 26 | 27 | 28 | 29 | 30 | 31 | 32 | 33 | 34 | 35 | 36 | 37 | 38 | 39 | 40 | 41 | 42 | 43 | 44 | 45 | 46 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         47 | 48 | 49 | 50 | 51 | 52 | 53 | 54 | 55 | 56 | 57 | 58 | 59 | 60 | 61 | 62 | 63 | 64 | 65 | 66 | 67 | 68 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *   

         69 | 70 | 71 | 72 | 73 | 74 | 75 | 76 | 77 | 78 | 79 | 80 | 81 | 82 | 83 | 84 | 85 | 86 | 87 | All
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|==1==
         *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *    *     *  

        Expression 89   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 90   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 91   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 92   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 93   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 94   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 95   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 96   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 97   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 98   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 99   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 100   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 101   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 102   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 103   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 104   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 105   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 106   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 107   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 108   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 109   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 110   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 111   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 112   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 113   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 114   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 115   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 116   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 117   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 118   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 119   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 120   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 121   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 122   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 123   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 124   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 125   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 126   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 127   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 128   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 129   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 130   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 131   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 132   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 133   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 134   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 135   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 136   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 137   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 138   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 139   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 140   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 141   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 142   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 143   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 144   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 145   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 146   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 147   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 148   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 149   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 150   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 151   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 152   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 153   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 154   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 155   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 156   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 157   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 158   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 159   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 160   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 161   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 162   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 163   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 164   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 165   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 166   (0/2)
        ^^^^^^^^^^^^^ - !=
         E | E
        =0=|=1=
         *   *

        Expression 167   (0/78)
        ^^^^^^^^^^^^^ - &&
         90 | 91 | 92 | 93 | 94 | 95 | 96 | 97 | 98 | 99 | 100 | 101 | 102 | 103 | 104 | 105 | 106 | 107 | 108 | 109 |
        =0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0==|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *    *    *    *    *    *    *    *    *    *    *     *     *     *     *     *     *     *     *     *    

         110 | 111 | 112 | 113 | 114 | 115 | 116 | 117 | 118 | 119 | 120 | 121 | 122 | 123 | 124 | 125 | 126 | 127 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         128 | 129 | 130 | 131 | 132 | 133 | 134 | 135 | 136 | 137 | 138 | 139 | 140 | 141 | 142 | 143 | 144 | 145 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         146 | 147 | 148 | 149 | 150 | 151 | 152 | 153 | 154 | 155 | 156 | 157 | 158 | 159 | 160 | 161 | 162 | 163 |
        =0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|=0===|
         *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *     *    

         164 | 165 | 166 | All
        =0===|=0===|=0===|==1==
         *     *     *      *  

        Expression 168   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 169   (0/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
