module main;

reg generate;

endmodule
