module main;

reg always_ff;

endmodule
