module main (
  a
);

input wire a;

endmodule
