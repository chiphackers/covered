module main;

parameter foo = 2 ** 3;

wire [(foo - 1):0] a;

endmodule
