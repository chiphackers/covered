module main #(parameter foo = 4); 

endmodule
