module dut_and( a, b, c );

output  a;
input   b;
input   c;

assign a = b & c;

endmodule
