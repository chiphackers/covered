module main;

reg always_comb;

endmodule
