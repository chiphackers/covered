module main;

reg bool;

endmodule
