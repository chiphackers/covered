/*
 Name:        timescale4.21.v
 Author:      Trevor Williams  (phase1geo@gmail.com)
 Date:        10/24/2008
 Purpose:     Verifies that real delays work properly when timescale is 10 s / 100 us
*/

`timescale 10 s / 100 us

module main;

reg a, b;

initial begin
	a = 1'b0;
	b = 1'b0;
	#(2.123_456_789_987_654);
	b = 1'b1;
	a = ($time == 64'd212346);
end

initial begin
`ifdef DUMP
        $dumpfile( "timescale4.21.vcd" );
        $dumpvars( 0, main );
`endif
        #(10);
        $finish;
end

endmodule
