module main;

reg        clk;
reg        reset;
reg        head1, head2;
reg        tail1, tail2;
reg        valid1, valid2;

fsma fsm1 (
  .clock( clk    ),
  .reset( reset  ),
  .head ( head1  ),
  .tail ( tail1  ),
  .valid( valid1 )
);

fsm fsm2 (
  .clock( clk    ),
  .reset( reset  ),
  .head ( head2  ),
  .tail ( tail2  ),
  .valid( valid2 )
);

initial begin
	$dumpfile( "fsm10.2.vcd" );
	$dumpvars( 0, main );
        reset  = 1'b1;
	head1  = 1'b0;
        tail1  = 1'b0;
        valid1 = 1'b0;
	head2  = 1'b0;
        tail2  = 1'b0;
        valid2 = 1'b0;
	#20;
	reset = 1'b0;
	#20;
	@(posedge clk);
        head1 <= 1'b1;
	valid1 <= 1'b1;
	@(posedge clk);
        head1 <= 1'b0;
	tail1 <= 1'b1;
	@(posedge clk);
	tail1  <= 1'b0;
	valid1 <= 1'b0;
	#20;
	$finish;
end

initial begin
	clk = 1'b0;
        forever #(2) clk = ~clk;
end

endmodule

/* HEADER
GROUPS fsm10.2 all iv vcd lxt
SIM    fsm10.2 all iv vcd  : iverilog -y ./lib fsm10.2.v; ./a.out                             : fsm10.2.vcd
SIM    fsm10.2 all iv lxt  : iverilog -y ./lib fsm10.2.v; ./a.out -lxt2; mv fsm10.2.vcd fsm10.2.lxt : fsm10.2.lxt
SCORE  fsm10.2.vcd     : -t main -vcd fsm10.2.vcd -o fsm10.2.cdd -y lib -v fsm10.2.v -F fsm=state,next_state : fsm10.2.cdd
SCORE  fsm10.2.lxt     : -t main -lxt fsm10.2.lxt -o fsm10.2.cdd -y lib -v fsm10.2.v -F fsm=state,next_state : fsm10.2.cdd
REPORT fsm10.2.cdd 1   : -d v -o fsm10.2.rptM fsm10.2.cdd                         : fsm10.2.rptM
REPORT fsm10.2.cdd 2   : -d v -w -o fsm10.2.rptWM fsm10.2.cdd                     : fsm10.2.rptWM
REPORT fsm10.2.cdd 3   : -d v -i -o fsm10.2.rptI fsm10.2.cdd                      : fsm10.2.rptI
REPORT fsm10.2.cdd 4   : -d v -w -i -o fsm10.2.rptWI fsm10.2.cdd                  : fsm10.2.rptWI
*/

/* OUTPUT fsm10.2.cdd
5 1 * 6 0 0 0 0
3 0 main main fsm10.2.v 1 56
2 1 52 7000a 1 0 20004 0 0 1 1 0
2 2 52 10003 0 1 400 0 0 clk
2 3 52 1000a 1 37 1006 1 2
2 4 53 1c001e 23 1 1c 0 0 clk
2 5 53 1b001b 23 1b 2002c 4 0 1 0 1102
2 6 53 150017 0 1 400 0 0 clk
2 7 53 15001e 23 37 602e 5 6
2 8 53 120012 1 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 9 53 120012 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 10 53 100013 47 2c 2000a 8 9 32 0 aa aa aa aa aa aa aa aa
1 clk 0 3 3000b 1 16 1102
1 reset 0 4 3000b 1 0 1002
1 head1 0 5 3000b 1 0 1102
1 head2 0 5 30012 1 0 2
1 tail1 0 6 3000b 1 0 1102
1 tail2 0 6 30012 1 0 2
1 valid1 0 7 3000b 1 0 1102
1 valid2 0 7 30013 1 0 2
4 7 10 10
4 10 7 0
4 3 10 10
3 0 fsma main.fsm1 lib/fsma.v 1 44
2 11 23 36003f 5 1 c 0 0 next_state
2 12 23 290032 1 32 4 0 0 #STATE_IDLE
2 13 23 210032 6 1a 200cc 11 12 32 0 33aa aa aa aa aa aa aa aa
2 14 23 210025 2 1 c 0 0 reset
2 15 23 21003f 6 19 201cc 13 14 2 0 330a
2 16 23 18001c 0 1 400 0 0 state
2 17 23 18003f 11 38 600e 15 16
2 18 23 110015 23 1 c 0 0 clock
2 19 23 9000f 0 2a 20000 0 0 2 0 a
2 20 23 90015 35 27 2100a 18 19 1 0 2
2 21 37 3d0046 1 32 4 0 0 #STATE_IDLE
2 22 37 300039 1 32 8 0 0 #STATE_HEAD
2 23 37 1f0039 3 1a 2010c 21 22 32 0 11aa aa aa aa aa aa aa aa
2 24 37 28002b 3 1 c 0 0 head
2 25 37 200024 3 1 c 0 0 valid
2 26 37 20002b 3 8 2024c 24 25 1 0 1102
2 27 37 1f0046 3 19 2024c 23 26 2 0 110a
2 28 37 12001b 0 1 400 0 0 next_state
2 29 37 120046 3 37 600e 27 28
2 30 38 3d0046 1 32 8 0 0 #STATE_DATA
2 31 38 300039 1 32 8 0 0 #STATE_TAIL
2 32 38 1f0039 1 1a 20208 30 31 32 0 aa aa aa aa aa aa aa aa
2 33 38 28002b 1 1 18 0 0 tail
2 34 38 200024 1 1 18 0 0 valid
2 35 38 20002b 1 8 20238 33 34 1 0 2
2 36 38 1f0046 1 19 20238 32 35 2 0 a
2 37 38 12001b 0 1 400 0 0 next_state
2 38 38 120046 1 37 602a 36 37
2 39 39 3d0046 0 32 10 0 0 #STATE_DATA
2 40 39 300039 0 32 10 0 0 #STATE_TAIL
2 41 39 1f0039 0 1a 20030 39 40 32 0 aa aa aa aa aa aa aa aa
2 42 39 28002b 0 1 10 0 0 tail
2 43 39 200024 0 1 10 0 0 valid
2 44 39 20002b 0 8 20030 42 43 1 0 2
2 45 39 1f0046 0 19 20030 41 44 2 0 a
2 46 39 12001b 0 1 400 0 0 next_state
2 47 39 120046 0 37 6022 45 46
2 48 40 3d0046 1 32 4 0 0 #STATE_IDLE
2 49 40 300039 1 32 8 0 0 #STATE_HEAD
2 50 40 1f0039 1 1a 20104 48 49 32 0 aa aa aa aa aa aa aa aa
2 51 40 28002b 1 1 4 0 0 head
2 52 40 200024 1 1 4 0 0 valid
2 53 40 20002b 1 8 20044 51 52 1 0 2
2 54 40 1f0046 1 19 20044 50 53 2 0 a
2 55 40 12001b 0 1 400 0 0 next_state
2 56 40 120046 1 37 6006 54 55
2 57 40 5000e 1 32 8 0 0 #STATE_TAIL
2 58 36 9000d d 1 e 0 0 state
2 59 40 0 2 2d 2420e 57 58 1 0 102
2 60 39 5000e 1 32 8 0 0 #STATE_DATA
2 61 39 0 2 2d 20206 60 58 1 0 2
2 62 38 5000e 1 32 8 0 0 #STATE_HEAD
2 63 38 0 3 2d 2020e 62 58 1 0 1102
2 64 37 5000e 1 32 4 0 0 #STATE_IDLE
2 65 37 0 6 2d 2014e 64 58 1 0 1102
2 66 34 230026 3 1 c 0 0 tail
2 67 34 230026 0 2a 20000 0 0 2 0 110a
2 68 34 230026 3 29 20008 66 67 1 0 2
2 69 34 1a001e 3 1 c 0 0 valid
2 70 34 1a001e 0 2a 20000 0 0 2 0 110a
2 71 34 1a001e 3 29 20008 69 70 1 0 2
2 72 34 120015 3 1 c 0 0 head
2 73 34 120015 0 2a 20000 0 0 2 0 110a
2 74 34 120015 3 29 20008 72 73 1 0 2
2 75 34 9000d 5 1 c 0 0 state
2 76 34 9000d 0 2a 20000 0 0 3 0 332a
2 77 34 9000d 5 29 20008 75 76 1 0 2
2 78 34 90015 6 2b 20008 74 77 1 0 2
2 79 34 9001e 6 2b 20008 71 78 1 0 2
2 80 34 90026 d 2b 2100a 68 79 1 0 2
2 81 0 0 5 1 f00e 0 0 next_state
2 82 0 0 5 1 f00e 0 0 state
1 #STATE_IDLE 0 0 0 32 0 0 0 0 0 0 0 0 0
1 #STATE_HEAD 0 0 0 32 0 1 0 0 0 0 0 0 0
1 #STATE_DATA 0 0 0 32 0 4 0 0 0 0 0 0 0
1 #STATE_TAIL 0 0 0 32 0 5 0 0 0 0 0 0 0
1 clock 0 9 a 1 0 1102
1 reset 0 10 a 1 0 1002
1 head 0 11 a 1 0 1102
1 tail 0 12 a 1 0 1102
1 valid 0 13 a 1 0 1102
1 state 0 20 3000b 2 0 330a
1 next_state 0 21 3000b 2 16 330a
4 82 82 82
4 81 81 81
4 17 20 20
4 20 17 0
4 56 80 80
4 59 56 80
4 47 80 80
4 61 47 59
4 38 80 80
4 63 38 61
4 29 80 80
4 65 29 63
4 80 65 0
6 82 81 1 02,08,08,0121,01,e1,c0,60014001a0018101
3 0 fsm main.fsm2 lib/fsm.v 1 35
2 83 23 36003f 1 1 4 0 0 next_state
2 84 23 290032 1 32 4 0 0 #STATE_IDLE
2 85 23 210032 2 1a 20044 83 84 32 0 aa aa aa aa aa aa aa aa
2 86 23 210025 2 1 c 0 0 reset
2 87 23 21003f 2 19 20144 85 86 2 0 a
2 88 23 18001c 0 1 400 0 0 state
2 89 23 18003f 11 38 6006 87 88
2 90 23 110015 23 1 c 0 0 clock
2 91 23 9000f 0 2a 20000 0 0 2 0 a
2 92 23 90015 35 27 2100a 90 91 1 0 2
2 93 28 3d0046 1 32 4 0 0 #STATE_IDLE
2 94 28 300039 1 32 8 0 0 #STATE_HEAD
2 95 28 1f0039 1 1a 20104 93 94 32 0 aa aa aa aa aa aa aa aa
2 96 28 28002b 1 1 4 0 0 head
2 97 28 200024 1 1 4 0 0 valid
2 98 28 20002b 1 8 20044 96 97 1 0 2
2 99 28 1f0046 1 19 20044 95 98 2 0 a
2 100 28 12001b 0 1 400 0 0 next_state
2 101 28 120046 1 37 6006 99 100
2 102 29 3d0046 0 32 10 0 0 #STATE_DATA
2 103 29 300039 0 32 10 0 0 #STATE_TAIL
2 104 29 1f0039 0 1a 20030 102 103 32 0 aa aa aa aa aa aa aa aa
2 105 29 28002b 0 1 10 0 0 tail
2 106 29 200024 0 1 10 0 0 valid
2 107 29 20002b 0 8 20030 105 106 1 0 2
2 108 29 1f0046 0 19 20030 104 107 2 0 a
2 109 29 12001b 0 1 400 0 0 next_state
2 110 29 120046 0 37 6022 108 109
2 111 30 3d0046 0 32 10 0 0 #STATE_DATA
2 112 30 300039 0 32 10 0 0 #STATE_TAIL
2 113 30 1f0039 0 1a 20030 111 112 32 0 aa aa aa aa aa aa aa aa
2 114 30 28002b 0 1 10 0 0 tail
2 115 30 200024 0 1 10 0 0 valid
2 116 30 20002b 0 8 20030 114 115 1 0 2
2 117 30 1f0046 0 19 20030 113 116 2 0 a
2 118 30 12001b 0 1 400 0 0 next_state
2 119 30 120046 0 37 6022 117 118
2 120 31 3d0046 0 32 10 0 0 #STATE_IDLE
2 121 31 300039 0 32 10 0 0 #STATE_HEAD
2 122 31 1f0039 0 1a 20030 120 121 32 0 aa aa aa aa aa aa aa aa
2 123 31 28002b 0 1 10 0 0 head
2 124 31 200024 0 1 10 0 0 valid
2 125 31 20002b 0 8 20030 123 124 1 0 2
2 126 31 1f0046 0 19 20030 122 125 2 0 a
2 127 31 12001b 0 1 400 0 0 next_state
2 128 31 120046 0 37 6022 126 127
2 129 31 5000e 1 32 8 0 0 #STATE_TAIL
2 130 27 9000d 5 1 6 0 0 state
2 131 31 0 1 2d 24006 129 130 1 0 2
2 132 30 5000e 1 32 8 0 0 #STATE_DATA
2 133 30 0 1 2d 20006 132 130 1 0 2
2 134 29 5000e 1 32 8 0 0 #STATE_HEAD
2 135 29 0 1 2d 20006 134 130 1 0 2
2 136 28 5000e 1 32 4 0 0 #STATE_IDLE
2 137 28 0 2 2d 2004e 136 130 1 0 102
2 138 25 230026 1 1 4 0 0 tail
2 139 25 230026 0 2a 20000 0 0 2 0 a
2 140 25 230026 1 29 20008 138 139 1 0 2
2 141 25 1a001e 1 1 4 0 0 valid
2 142 25 1a001e 0 2a 20000 0 0 2 0 a
2 143 25 1a001e 1 29 20008 141 142 1 0 2
2 144 25 120015 1 1 4 0 0 head
2 145 25 120015 0 2a 20000 0 0 2 0 a
2 146 25 120015 1 29 20008 144 145 1 0 2
2 147 25 9000d 2 1 4 0 0 state
2 148 25 9000d 0 2a 20000 0 0 3 0 2a
2 149 25 9000d 2 29 20008 147 148 1 0 2
2 150 25 90015 2 2b 20008 146 149 1 0 2
2 151 25 9001e 2 2b 20008 143 150 1 0 2
2 152 25 90026 5 2b 2100a 140 151 1 0 2
2 153 0 0 1 1 f006 0 0 next_state
2 154 0 0 2 1 f006 0 0 state
1 #STATE_IDLE 0 0 0 32 0 0 0 0 0 0 0 0 0
1 #STATE_HEAD 0 0 0 32 0 1 0 0 0 0 0 0 0
1 #STATE_DATA 0 0 0 32 0 4 0 0 0 0 0 0 0
1 #STATE_TAIL 0 0 0 32 0 5 0 0 0 0 0 0 0
1 clock 0 9 a 1 0 1102
1 reset 0 10 a 1 0 1002
1 head 0 11 a 1 0 2
1 tail 0 12 a 1 0 2
1 valid 0 13 a 1 0 2
1 state 0 20 3000b 2 0 a
1 next_state 0 21 3000b 2 16 a
4 154 154 154
4 153 153 153
4 89 92 92
4 92 89 0
4 128 152 152
4 131 128 152
4 119 152 152
4 133 119 131
4 110 152 152
4 135 110 133
4 101 152 152
4 137 101 135
4 152 137 0
6 154 153 1 02,02,01,,01,
*/

/* OUTPUT fsm10.2.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm10.2.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm10.2.v                  2/    0/    2      100%
  fsma                    fsma.v                     6/    1/    7       86%
  fsm                     fsm.v                      4/    3/    7       57%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           39:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA


    Module: fsm, File: lib/fsm.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           29:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
           30:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
           31:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm10.2.v                  4/    4/    8       50%             5/    3/    8       62%
  fsma                    fsma.v                     8/    1/    9       89%             9/    0/    9      100%
  fsm                     fsm.v                      1/    8/    9       11%             2/    7/    9       22%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm10.2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      head2                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      tail2                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      valid2                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: fsma, File: lib/fsma.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: fsm, File: lib/fsm.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      head                      0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      tail                      0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      valid                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      state                     0->1: 2'h0
      ......................... 1->0: 2'h0 ...
      next_state                0->1: 2'h0
      ......................... 1->0: 2'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm10.2.v                           2/   0/   2      100%
  fsma                              fsma.v                             19/  16/  35       54%
  fsm                               fsm.v                              11/  24/  35       31%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             37:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             38:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             39:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             40:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *


    Module: fsm, File: lib/fsm.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    state <= reset ? STATE_IDLE : next_state
                             |--------------1--------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    case( state ) 
                          |-1-|   
                    STATE_IDLE :

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             30:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm10.2.v                 0/   0/   0      100%            0/   0/   0      100%
  fsma                    fsma.v                    3/   1/   4       75%            4/   4/   8       50%
  fsm                     fsm.v                     1/  ? /  ?        ? %            1/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          2'h2

        Missed State Transitions

          From State    To State  
          ==========    ==========
          2'h1       -> 2'h2      
          2'h2       -> 2'h3      
          2'h2       -> 2'h2      
          2'h3       -> 2'h1      


    Module: fsm, File: lib/fsm.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          2'h0

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      



*/

/* OUTPUT fsm10.2.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm10.2.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm10.2.v                  2/    0/    2      100%
  fsma                    fsma.v                     6/    1/    7       86%
  fsm                     fsm.v                      4/    3/    7       57%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           39:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA


    Module: fsm, File: lib/fsm.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           29:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
           30:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
           31:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm10.2.v                  4/    4/    8       50%             5/    3/    8       62%
  fsma                    fsma.v                     8/    1/    9       89%             9/    0/    9      100%
  fsm                     fsm.v                      1/    8/    9       11%             2/    7/    9       22%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm10.2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      head2                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      tail2                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      valid2                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: fsma, File: lib/fsma.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: fsm, File: lib/fsm.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      head                      0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      tail                      0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      valid                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      state                     0->1: 2'h0
      ......................... 1->0: 2'h0 ...
      next_state                0->1: 2'h0
      ......................... 1->0: 2'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm10.2.v                           2/   0/   2      100%
  fsma                              fsma.v                             19/  16/  35       54%
  fsm                               fsm.v                              11/  24/  35       31%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             37:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             38:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             39:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             40:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *


    Module: fsm, File: lib/fsm.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    state <= reset ? STATE_IDLE : next_state
                             |--------------1--------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    case( state ) STATE_IDLE :
                          |-1-|               

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             30:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm10.2.v                 0/   0/   0      100%            0/   0/   0      100%
  fsma                    fsma.v                    3/   1/   4       75%            4/   4/   8       50%
  fsm                     fsm.v                     1/  ? /  ?        ? %            1/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          2'h2

        Missed State Transitions

          From State    To State  
          ==========    ==========
          2'h1       -> 2'h2      
          2'h2       -> 2'h3      
          2'h2       -> 2'h2      
          2'h3       -> 2'h1      


    Module: fsm, File: lib/fsm.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          2'h0

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      



*/

/* OUTPUT fsm10.2.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm10.2.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          2/    0/    2      100%
  <NA>.main.fsm1                                     6/    1/    7       86%
  <NA>.main.fsm2                                     4/    3/    7       57%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           39:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA


    Module: fsm, File: lib/fsm.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           29:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
           30:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
           31:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          4/    4/    8       50%             5/    3/    8       62%
  <NA>.main.fsm1                                     8/    1/    9       89%             9/    0/    9      100%
  <NA>.main.fsm2                                     1/    8/    9       11%             2/    7/    9       22%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm10.2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      head2                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      tail2                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      valid2                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: fsma, File: lib/fsma.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: fsm, File: lib/fsm.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      head                      0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      tail                      0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      valid                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      state                     0->1: 2'h0
      ......................... 1->0: 2'h0 ...
      next_state                0->1: 2'h0
      ......................... 1->0: 2'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             2/   0/   2      100%
  <NA>.main.fsm1                                                       19/  16/  35       54%
  <NA>.main.fsm2                                                       11/  24/  35       31%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             37:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             38:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             39:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             40:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *


    Module: fsm, File: lib/fsm.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    state <= reset ? STATE_IDLE : next_state
                             |--------------1--------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    case( state ) 
                          |-1-|   
                    STATE_IDLE :

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             30:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.fsm1                                    3/   1/   4       75%            4/   4/   8       50%
  <NA>.main.fsm2                                    1/  ? /  ?        ? %            1/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          2'h2

        Missed State Transitions

          From State    To State  
          ==========    ==========
          2'h1       -> 2'h2      
          2'h2       -> 2'h3      
          2'h2       -> 2'h2      
          2'h3       -> 2'h1      


    Module: fsm, File: lib/fsm.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          2'h0

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      



*/

/* OUTPUT fsm10.2.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm10.2.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          2/    0/    2      100%
  <NA>.main.fsm1                                     6/    1/    7       86%
  <NA>.main.fsm2                                     4/    3/    7       57%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           39:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA


    Module: fsm, File: lib/fsm.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           29:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
           30:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
           31:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          4/    4/    8       50%             5/    3/    8       62%
  <NA>.main.fsm1                                     8/    1/    9       89%             9/    0/    9      100%
  <NA>.main.fsm2                                     1/    8/    9       11%             2/    7/    9       22%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm10.2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      head2                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      tail2                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      valid2                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: fsma, File: lib/fsma.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: fsm, File: lib/fsm.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      head                      0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      tail                      0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      valid                     0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      state                     0->1: 2'h0
      ......................... 1->0: 2'h0 ...
      next_state                0->1: 2'h0
      ......................... 1->0: 2'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             2/   0/   2      100%
  <NA>.main.fsm1                                                       19/  16/  35       54%
  <NA>.main.fsm2                                                       11/  24/  35       31%
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             37:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             38:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             39:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             40:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *


    Module: fsm, File: lib/fsm.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    state <= reset ? STATE_IDLE : next_state
                             |--------------1--------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    case( state ) STATE_IDLE :
                          |-1-|               

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             30:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.fsm1                                    3/   1/   4       75%            4/   4/   8       50%
  <NA>.main.fsm2                                    1/  ? /  ?        ? %            1/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: fsma, File: lib/fsma.v, Instance: <NA>.main.fsm1
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Missed States

          States
          ======
          2'h2

        Missed State Transitions

          From State    To State  
          ==========    ==========
          2'h1       -> 2'h2      
          2'h2       -> 2'h3      
          2'h2       -> 2'h2      
          2'h3       -> 2'h1      


    Module: fsm, File: lib/fsm.v, Instance: <NA>.main.fsm2
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          2'h0

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      



*/
