module main;

wire a;

always_comb
  $display( "HERE!" );
	  
/*
initial begin
	#10;
	$finish;
end
*/

endmodule
