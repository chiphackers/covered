module main;

reg a, b;

initial begin : foobar
	a = 1'b0;
end

initial begin : barfoo
	b <= 1'b1;
end

initial begin
	#10;
	begin : fooey
	 reg c, d;
	 c <= a & b;
	 d <= a | b;
	end
	begin : barry
         reg e, f;
	 e <= a ^ b;
	 f <= a ~^ b;
	end
end

initial begin
        $dumpfile( "named_block1.vcd" );
        $dumpvars( 0, main );
        #100;
        $finish;
end

endmodule

/* HEADER
GROUPS named_block1 all iv vcs vcd lxt
SIM    named_block1 all iv vcd  : iverilog named_block1.v; ./a.out                             : named_block1.vcd
SIM    named_block1 all iv lxt  : iverilog named_block1.v; ./a.out -lxt2; mv named_block1.vcd named_block1.lxt : named_block1.lxt
SIM    named_block1 all vcs vcd : vcs named_block1.v; ./simv                                   : named_block1.vcd
SCORE  named_block1.vcd     : -t main -vcd named_block1.vcd -o named_block1.cdd -v named_block1.v : named_block1.cdd
SCORE  named_block1.lxt     : -t main -lxt named_block1.lxt -o named_block1.cdd -v named_block1.v : named_block1.cdd
REPORT named_block1.cdd 1   : -d v -o named_block1.rptM named_block1.cdd                         : named_block1.rptM
REPORT named_block1.cdd 2   : -d v -w -o named_block1.rptWM named_block1.cdd                     : named_block1.rptWM
REPORT named_block1.cdd 3   : -d v -i -o named_block1.rptI named_block1.cdd                      : named_block1.rptI
REPORT named_block1.cdd 4   : -d v -w -i -o named_block1.rptWI named_block1.cdd                  : named_block1.rptWI
*/

/* OUTPUT named_block1.cdd
5 1 * 6 0 0 0 0
3 0 main main named_block1.v 1 34
2 1 5 8000c 2 3d 2100a 0 0 1 0 2 foobar
2 2 9 8000c 2 3d 2100a 0 0 1 0 2 barfoo
2 3 14 20003 1 0 20008 0 0 32 64 44 0 0 0 0 0 0 0
2 4 14 20003 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 5 14 10003 2 2c 2100a 3 4 32 0 aa aa aa aa aa aa aa aa
2 6 15 10005 2 3d 2000a 0 0 1 0 2 fooey
2 7 20 10005 2 3d 2000a 0 0 1 0 2 barry
1 a 0 3 30004 1 16 2
1 b 0 3 30007 1 0 2
4 1 0 0
4 2 0 0
4 7 0 0
4 6 7 0
4 5 6 0
3 1 main.foobar main.foobar named_block1.v 5 7
2 8 6 50008 1 0 20004 0 0 1 1 0
2 9 6 10001 0 1 400 0 0 a
2 10 6 10008 1 37 11006 8 9
4 10 0 0
3 1 main.barfoo main.barfoo named_block1.v 9 11
2 11 10 60009 1 0 20008 0 0 1 1 1
2 12 10 10001 0 1 400 0 0 b
2 13 10 10009 1 38 1100a 11 12
4 13 0 0
3 1 main.fooey main.fooey named_block1.v 15 19
2 14 17 b000b 1 1 8 0 0 b
2 15 17 70007 1 1 4 0 0 a
2 16 17 7000b 1 8 20084 14 15 1 0 2
2 17 17 20002 0 1 400 0 0 c
2 18 17 2000b 1 38 11006 16 17
2 19 18 b000b 1 1 8 0 0 b
2 20 18 70007 1 1 4 0 0 a
2 21 18 7000b 1 9 20088 19 20 1 0 2
2 22 18 20002 0 1 400 0 0 d
2 23 18 2000b 1 38 a 21 22
1 c 0 16 30006 1 0 2
1 d 0 16 30009 1 0 2
4 23 0 0
4 18 23 23
3 1 main.barry main.barry named_block1.v 20 24
2 24 22 b000b 1 1 8 0 0 b
2 25 22 70007 1 1 4 0 0 a
2 26 22 7000b 1 2 20088 24 25 1 0 2
2 27 22 20002 0 1 400 0 0 e
2 28 22 2000b 1 38 1100a 26 27
2 29 23 c000c 1 1 8 0 0 b
2 30 23 70007 1 1 4 0 0 a
2 31 23 7000c 1 c 20084 29 30 1 0 2
2 32 23 20002 0 1 400 0 0 f
2 33 23 2000c 1 38 6 31 32
1 e 0 21 3000d 1 0 2
1 f 0 21 30010 1 0 2
4 33 0 0
4 28 33 33
*/

/* OUTPUT named_block1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : named_block1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    named_block1.v             0/    0/    0      100%
  main.foobar             named_block1.v             1/    0/    1      100%
  main.barfoo             named_block1.v             1/    0/    1      100%
  main.fooey              named_block1.v             2/    0/    2      100%
  main.barry              named_block1.v             2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    named_block1.v             0/    2/    2        0%             0/    2/    2        0%
  main.foobar             named_block1.v             0/    0/    0      100%             0/    0/    0      100%
  main.barfoo             named_block1.v             0/    0/    0      100%             0/    0/    0      100%
  main.fooey              named_block1.v             0/    2/    2        0%             0/    2/    2        0%
  main.barry              named_block1.v             0/    2/    2        0%             0/    2/    2        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Named Block: main.fooey, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Named Block: main.barry, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              named_block1.v                      0/   0/   0      100%
  main.foobar                       named_block1.v                      0/   0/   0      100%
  main.barfoo                       named_block1.v                      0/   0/   0      100%
  main.fooey                        named_block1.v                      2/   6/   8       25%
  main.barry                        named_block1.v                      2/   6/   8       25%
---------------------------------------------------------------------------------------------------------------------

    Named Block: main.fooey, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             17:     c  <= ( a  &  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             18:     d  <= ( a  |  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *


    Named Block: main.barry, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:     e  <= ( a  ^  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:     f  <= ( a  ~^  b )
                           |----1-----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ~^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    named_block1.v            0/   0/   0      100%            0/   0/   0      100%
  main.foobar             named_block1.v            0/   0/   0      100%            0/   0/   0      100%
  main.barfoo             named_block1.v            0/   0/   0      100%            0/   0/   0      100%
  main.fooey              named_block1.v            0/   0/   0      100%            0/   0/   0      100%
  main.barry              named_block1.v            0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT named_block1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : named_block1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    named_block1.v             0/    0/    0      100%
  main.foobar             named_block1.v             1/    0/    1      100%
  main.barfoo             named_block1.v             1/    0/    1      100%
  main.fooey              named_block1.v             2/    0/    2      100%
  main.barry              named_block1.v             2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    named_block1.v             0/    2/    2        0%             0/    2/    2        0%
  main.foobar             named_block1.v             0/    0/    0      100%             0/    0/    0      100%
  main.barfoo             named_block1.v             0/    0/    0      100%             0/    0/    0      100%
  main.fooey              named_block1.v             0/    2/    2        0%             0/    2/    2        0%
  main.barry              named_block1.v             0/    2/    2        0%             0/    2/    2        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Named Block: main.fooey, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Named Block: main.barry, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              named_block1.v                      0/   0/   0      100%
  main.foobar                       named_block1.v                      0/   0/   0      100%
  main.barfoo                       named_block1.v                      0/   0/   0      100%
  main.fooey                        named_block1.v                      2/   6/   8       25%
  main.barry                        named_block1.v                      2/   6/   8       25%
---------------------------------------------------------------------------------------------------------------------

    Named Block: main.fooey, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             17:     c  <= ( a  &  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             18:     d  <= ( a  |  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *


    Named Block: main.barry, File: named_block1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:     e  <= ( a  ^  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:     f  <= ( a  ~^  b )
                           |----1-----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ~^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    named_block1.v            0/   0/   0      100%            0/   0/   0      100%
  main.foobar             named_block1.v            0/   0/   0      100%            0/   0/   0      100%
  main.barfoo             named_block1.v            0/   0/   0      100%            0/   0/   0      100%
  main.fooey              named_block1.v            0/   0/   0      100%            0/   0/   0      100%
  main.barry              named_block1.v            0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT named_block1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : named_block1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%
  <NA>.main.foobar                                   1/    0/    1      100%
  <NA>.main.barfoo                                   1/    0/    1      100%
  <NA>.main.fooey                                    2/    0/    2      100%
  <NA>.main.barry                                    2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.foobar                                   0/    0/    0      100%             0/    0/    0      100%
  <NA>.main.barfoo                                   0/    0/    0      100%             0/    0/    0      100%
  <NA>.main.fooey                                    0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.barry                                    0/    2/    2        0%             0/    2/    2        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: named_block1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Named Block: main.fooey, File: named_block1.v, Instance: <NA>.main.fooey
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Named Block: main.barry, File: named_block1.v, Instance: <NA>.main.barry
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%
  <NA>.main.foobar                                                      0/   0/   0      100%
  <NA>.main.barfoo                                                      0/   0/   0      100%
  <NA>.main.fooey                                                       2/   6/   8       25%
  <NA>.main.barry                                                       2/   6/   8       25%
---------------------------------------------------------------------------------------------------------------------

    Named Block: main.fooey, File: named_block1.v, Instance: <NA>.main.fooey
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             17:     c  <= ( a  &  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             18:     d  <= ( a  |  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *


    Named Block: main.barry, File: named_block1.v, Instance: <NA>.main.barry
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:     e  <= ( a  ^  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:     f  <= ( a  ~^  b )
                           |----1-----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ~^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.foobar                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.barfoo                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.fooey                                   0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.barry                                   0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT named_block1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : named_block1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%
  <NA>.main.foobar                                   1/    0/    1      100%
  <NA>.main.barfoo                                   1/    0/    1      100%
  <NA>.main.fooey                                    2/    0/    2      100%
  <NA>.main.barry                                    2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.foobar                                   0/    0/    0      100%             0/    0/    0      100%
  <NA>.main.barfoo                                   0/    0/    0      100%             0/    0/    0      100%
  <NA>.main.fooey                                    0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.barry                                    0/    2/    2        0%             0/    2/    2        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: named_block1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Named Block: main.fooey, File: named_block1.v, Instance: <NA>.main.fooey
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Named Block: main.barry, File: named_block1.v, Instance: <NA>.main.barry
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      e                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%
  <NA>.main.foobar                                                      0/   0/   0      100%
  <NA>.main.barfoo                                                      0/   0/   0      100%
  <NA>.main.fooey                                                       2/   6/   8       25%
  <NA>.main.barry                                                       2/   6/   8       25%
---------------------------------------------------------------------------------------------------------------------

    Named Block: main.fooey, File: named_block1.v, Instance: <NA>.main.fooey
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             17:     c  <= ( a  &  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             18:     d  <= ( a  |  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - |
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *


    Named Block: main.barry, File: named_block1.v, Instance: <NA>.main.barry
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:     e  <= ( a  ^  b )
                           |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:     f  <= ( a  ~^  b )
                           |----1-----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ~^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *         *    *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.foobar                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.barfoo                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.fooey                                   0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.barry                                   0/   0/   0      100%            0/   0/   0      100%


*/
