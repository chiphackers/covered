module main (
  a
);

output reg a;

endmodule
