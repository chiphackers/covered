module main;

foo bar[3:0]();

endmodule

//------------------------

module foo;

wire a;

endmodule
