module main;

parameter STATE_IDLE = 2'b00,
          STATE_HEAD = 2'b01,
          STATE_DATA = 2'b10,
          STATE_TAIL = 2'b11;

reg        clk;
reg        reset;
reg        head;
reg        tail;
reg        valid;
reg [1:0]  state;
reg [1:0]  next_state;

always @(posedge clk) state <= reset ? STATE_IDLE : next_state;

(* covered_fsm, channel, is="state", os="next_state",
                         trans="STATE_IDLE->STATE_HEAD",
                         trans="STATE_IDLE->STATE_IDLE" *)
always @(state or head or valid or tail)
  begin
   case( state )
     STATE_IDLE:  next_state = (valid & head) ? STATE_HEAD : STATE_IDLE;
     STATE_HEAD:  next_state = (valid & tail) ? STATE_TAIL : STATE_DATA;
     STATE_DATA:  next_state = (valid & tail) ? STATE_TAIL : STATE_DATA;
     STATE_TAIL:  next_state = (valid & head) ? STATE_HEAD : STATE_IDLE;
   endcase
  end

initial begin
	$dumpfile( "fsm7.4.vcd" );
	$dumpvars( 0, main );
        reset = 1'b1;
	head  = 1'b0;
        tail  = 1'b0;
        valid = 1'b0;
	#20;
	reset = 1'b0;
	#20;
	@(posedge clk);
        head <= 1'b1;
	valid <= 1'b1;
	@(posedge clk);
        head <= 1'b0;
	tail <= 1'b1;
	@(posedge clk);
	tail  <= 1'b0;
	valid <= 1'b0;
	#20;
	$finish;
end

initial begin
	clk = 1'b0;
        forever #(2) clk = ~clk;
end

endmodule

/* HEADER
GROUPS fsm7.4 all iv vcd lxt
SIM    fsm7.4 all iv vcd  : iverilog fsm7.4.v; ./a.out                             : fsm7.4.vcd
SIM    fsm7.4 all iv lxt  : iverilog fsm7.4.v; ./a.out -lxt2; mv fsm7.4.vcd fsm7.4.lxt : fsm7.4.lxt
SCORE  fsm7.4.vcd     : -t main -vcd fsm7.4.vcd -o fsm7.4.cdd -v fsm7.4.v : fsm7.4.cdd
SCORE  fsm7.4.lxt     : -t main -lxt fsm7.4.lxt -o fsm7.4.cdd -v fsm7.4.v : fsm7.4.cdd
REPORT fsm7.4.cdd 1   : -d v -o fsm7.4.rptM fsm7.4.cdd                         : fsm7.4.rptM
REPORT fsm7.4.cdd 2   : -d v -w -o fsm7.4.rptWM fsm7.4.cdd                     : fsm7.4.rptWM
REPORT fsm7.4.cdd 3   : -d v -i -o fsm7.4.rptI fsm7.4.cdd                      : fsm7.4.rptI
REPORT fsm7.4.cdd 4   : -d v -w -i -o fsm7.4.rptWI fsm7.4.cdd                  : fsm7.4.rptWI
*/

/* OUTPUT fsm7.4.cdd
5 1 * 6 0 0 0 0
3 0 main main fsm7.4.v 1 59
2 1 16 34003d 5 1 c 0 0 next_state
2 2 16 270030 1 32 4 0 0 #STATE_IDLE
2 3 16 1f0030 7 1a 200cc 1 2 32 0 33aa aa aa aa aa aa aa aa
2 4 16 1f0023 2 1 c 0 0 reset
2 5 16 1f003d 7 19 201cc 3 4 2 0 330a
2 6 16 16001a 0 1 400 0 0 state
2 7 16 16003d 12 38 600e 5 6
2 8 16 110013 24 1 c 0 0 clk
2 9 16 9000f 0 2a 20000 0 0 2 0 a
2 10 16 90013 37 27 2100a 8 9 1 0 2
2 11 24 3d0046 1 32 4 0 0 #STATE_IDLE
2 12 24 300039 1 32 8 0 0 #STATE_HEAD
2 13 24 1f0039 3 1a 2010c 11 12 32 0 11aa aa aa aa aa aa aa aa
2 14 24 28002b 3 1 c 0 0 head
2 15 24 200024 3 1 c 0 0 valid
2 16 24 20002b 3 8 2024c 14 15 1 0 1102
2 17 24 1f0046 3 19 2024c 13 16 2 0 110a
2 18 24 12001b 0 1 400 0 0 next_state
2 19 24 120046 3 37 600e 17 18
2 20 25 3d0046 1 32 8 0 0 #STATE_DATA
2 21 25 300039 1 32 8 0 0 #STATE_TAIL
2 22 25 1f0039 1 1a 20208 20 21 32 0 aa aa aa aa aa aa aa aa
2 23 25 28002b 1 1 18 0 0 tail
2 24 25 200024 1 1 18 0 0 valid
2 25 25 20002b 1 8 20238 23 24 1 0 2
2 26 25 1f0046 1 19 20238 22 25 2 0 a
2 27 25 12001b 0 1 400 0 0 next_state
2 28 25 120046 1 37 602a 26 27
2 29 26 3d0046 0 32 10 0 0 #STATE_DATA
2 30 26 300039 0 32 10 0 0 #STATE_TAIL
2 31 26 1f0039 0 1a 20030 29 30 32 0 aa aa aa aa aa aa aa aa
2 32 26 28002b 0 1 10 0 0 tail
2 33 26 200024 0 1 10 0 0 valid
2 34 26 20002b 0 8 20030 32 33 1 0 2
2 35 26 1f0046 0 19 20030 31 34 2 0 a
2 36 26 12001b 0 1 400 0 0 next_state
2 37 26 120046 0 37 6022 35 36
2 38 27 3d0046 1 32 4 0 0 #STATE_IDLE
2 39 27 300039 1 32 8 0 0 #STATE_HEAD
2 40 27 1f0039 1 1a 20104 38 39 32 0 aa aa aa aa aa aa aa aa
2 41 27 28002b 1 1 4 0 0 head
2 42 27 200024 1 1 4 0 0 valid
2 43 27 20002b 1 8 20044 41 42 1 0 2
2 44 27 1f0046 1 19 20044 40 43 2 0 a
2 45 27 12001b 0 1 400 0 0 next_state
2 46 27 120046 1 37 6006 44 45
2 47 27 5000e 1 32 8 0 0 #STATE_TAIL
2 48 23 9000d d 1 e 0 0 state
2 49 27 0 2 2d 2420e 47 48 1 0 102
2 50 26 5000e 1 32 8 0 0 #STATE_DATA
2 51 26 0 2 2d 20206 50 48 1 0 2
2 52 25 5000e 1 32 8 0 0 #STATE_HEAD
2 53 25 0 3 2d 2020e 52 48 1 0 1102
2 54 24 5000e 1 32 4 0 0 #STATE_IDLE
2 55 24 0 6 2d 2014e 54 48 1 0 1102
2 56 21 230026 3 1 c 0 0 tail
2 57 21 230026 0 2a 20000 0 0 2 0 110a
2 58 21 230026 3 29 20008 56 57 1 0 2
2 59 21 1a001e 3 1 c 0 0 valid
2 60 21 1a001e 0 2a 20000 0 0 2 0 110a
2 61 21 1a001e 3 29 20008 59 60 1 0 2
2 62 21 120015 3 1 c 0 0 head
2 63 21 120015 0 2a 20000 0 0 2 0 110a
2 64 21 120015 3 29 20008 62 63 1 0 2
2 65 21 9000d 5 1 c 0 0 state
2 66 21 9000d 0 2a 20000 0 0 3 0 332a
2 67 21 9000d 5 29 20008 65 66 1 0 2
2 68 21 90015 6 2b 20008 64 67 1 0 2
2 69 21 9001e 6 2b 20008 61 68 1 0 2
2 70 21 90026 d 2b 2100a 58 69 1 0 2
2 71 55 7000a 1 0 20004 0 0 1 1 0
2 72 55 10003 0 1 400 0 0 clk
2 73 55 1000a 1 37 1006 71 72
2 74 56 1c001e 23 1 1c 0 0 clk
2 75 56 1b001b 23 1b 2002c 74 0 1 0 1102
2 76 56 150017 0 1 400 0 0 clk
2 77 56 15001e 23 37 602e 75 76
2 78 56 120012 1 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 79 56 120012 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 80 56 100013 47 2c 2000a 78 79 32 0 aa aa aa aa aa aa aa aa
2 81 0 0 5 1 f00e 0 0 next_state
2 82 0 0 5 1 f00e 0 0 state
1 #STATE_IDLE 0 0 0 32 0 0 0 0 0 0 0 0 0
1 #STATE_HEAD 0 0 0 32 0 1 0 0 0 0 0 0 0
1 #STATE_DATA 0 0 0 32 0 4 0 0 0 0 0 0 0
1 #STATE_TAIL 0 0 0 32 0 5 0 0 0 0 0 0 0
1 clk 0 8 3000b 1 16 1102
1 reset 0 9 3000b 1 0 1002
1 head 0 10 3000b 1 0 1102
1 tail 0 11 3000b 1 0 1102
1 valid 0 12 3000b 1 0 1102
1 state 0 13 3000b 2 0 330a
1 next_state 0 14 3000b 2 16 330a
4 82 82 82
4 81 81 81
4 7 10 10
4 10 7 0
4 46 70 70
4 49 46 70
4 37 70 70
4 51 37 49
4 28 70 70
4 53 28 51
4 19 70 70
4 55 19 53
4 70 55 0
4 77 80 80
4 80 77 0
4 73 80 80
6 82 81 1 02,04,04,0121,01,e1,8101
*/

/* OUTPUT fsm7.4.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm7.4.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.4.v                   8/    1/    9       89%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           26:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.4.v                   8/    1/    9       89%             9/    0/    9      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm7.4.v                           21/  16/  37       57%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.4.v                  3/   0/   3      100%            4/   0/   4      100%


*/

/* OUTPUT fsm7.4.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm7.4.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.4.v                   8/    1/    9       89%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           26:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.4.v                   8/    1/    9       89%             9/    0/    9      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm7.4.v                           21/  16/  37       57%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm7.4.v                  3/   0/   3      100%            4/   0/   4      100%


*/

/* OUTPUT fsm7.4.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm7.4.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          8/    1/    9       89%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           26:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          8/    1/    9       89%             9/    0/    9      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            21/  16/  37       57%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         3/   0/   3      100%            4/   0/   4      100%


*/

/* OUTPUT fsm7.4.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm7.4.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          8/    1/    9       89%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           26:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          8/    1/    9       89%             9/    0/    9      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            21/  16/  37       57%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm7.4.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         3/   0/   3      100%            4/   0/   4      100%


*/
