module main;

reg [31:0] a;
reg        b;

initial begin
        a = 0;
        b = 1'b0;
	do
          begin
           #5;
           if( !a[1] )
             a = a + 2;
           else
             a = a + 1;
          end
        while( a < 10 );
	b = 1'b1;
end

initial begin
        $dumpfile( "do_while1.vcd" );
        $dumpvars( 0, main );
        #20;
        $finish;
end

endmodule
