module level3b(
  input  wire a,
  output wire b
);

assign b = ~a;

endmodule
