module main;

reg	[3:0]	a;
reg	[3:0]	b;
wire	[3:0]	z;
wire		carry;
wire	[4:0]	result;

assign result = {carry, z};

adder4 add( a, b, carry, z );

initial begin
	$dumpfile( "instance2.vcd" );
	$dumpvars( 0, main );
	a = 4'h0;
	b = 4'h1;
	#5;
	a = 4'h8;
	b = 4'h4;
	#5;
	b = 4'h8;
	#5;
	$finish;
end

endmodule

/* HEADER
GROUPS instance2 all iv vcs vcd lxt
SIM    instance2 all iv vcd  : iverilog -y ./lib instance2.v; ./a.out                             : instance2.vcd
SIM    instance2 all iv lxt  : iverilog -y ./lib instance2.v; ./a.out -lxt2; mv instance2.vcd instance2.lxt : instance2.lxt
SIM    instance2 all vcs vcd : vcs +libext+.v+ -y ./lib instance2.v; ./simv                                 : instance2.vcd
SCORE  instance2.vcd     : -t main -vcd instance2.vcd -o instance2.cdd -v instance2.v -y ./lib : instance2.cdd
SCORE  instance2.lxt     : -t main -lxt instance2.lxt -o instance2.cdd -v instance2.v -y ./lib : instance2.cdd
REPORT instance2.cdd 1   : -d v -o instance2.rptM instance2.cdd                         : instance2.rptM
REPORT instance2.cdd 2   : -d v -w -o instance2.rptWM instance2.cdd                     : instance2.rptWM
REPORT instance2.cdd 3   : -d v -i -o instance2.rptI instance2.cdd                      : instance2.rptI
REPORT instance2.cdd 4   : -d v -w -i -o instance2.rptWI instance2.cdd                  : instance2.rptWI
*/

/* OUTPUT instance2.cdd
5 1 * 6 0 0 0 0
3 0 main main instance2.v 1 27
2 1 9 180018 3 1 c 0 0 z
2 2 9 110015 2 1 c 0 0 carry
2 3 9 110018 3 31 20188 1 2 5 0 dcaa 102
2 4 9 100019 3 26 20008 3 0 5 0 dcaa 102
2 5 9 7000c 0 1 400 0 0 result
2 6 9 70019 3 35 f00a 4 5
1 a 0 3 3000a 4 0 8aa
1 b 0 4 3000a 4 0 5caa
1 z 0 5 3000b 4 0 dcaa
1 carry 0 6 30006 1 0 102
1 result 0 7 3000b 5 0 dcaa 102
4 6 6 6
3 0 adder4 main.add ./lib/adder4.v 1 22
1 a 0 8 c 4 0 8aa
1 b 0 9 c 4 0 5caa
1 c 0 10 10008 1 0 102
1 z 0 11 1000f 4 0 dcaa
1 c0 0 13 30009 1 0 2
1 c1 0 13 3000d 1 0 2
1 c2 0 13 30011 1 0 2
3 0 adder1 main.add.bit0 ./lib/adder1.v 1 18
2 7 15 f000f 2 1 c 0 0 b
2 8 15 b000b 1 1 4 0 0 a
2 9 15 b000f 2 2 200cc 7 8 1 0 1002
2 10 15 70007 0 1 400 0 0 z
2 11 15 7000f 2 35 f00e 9 10
2 12 16 f000f 2 1 c 0 0 b
2 13 16 b000b 1 1 4 0 0 a
2 14 16 b000f 2 8 200c4 12 13 1 0 2
2 15 16 70007 0 1 400 0 0 c
2 16 16 7000f 1 35 f006 14 15
1 a 0 8 7 1 0 2
1 b 0 9 7 1 0 1002
1 c 0 10 10008 1 0 2
1 z 0 11 10009 1 0 1002
4 11 11 11
4 16 16 16
3 0 adder1 main.add.bit1 ./lib/adder1.v 1 18
2 17 15 f000f 1 1 4 0 0 b
2 18 15 b000b 1 1 4 0 0 a
2 19 15 b000f 1 2 20044 17 18 1 0 2
2 20 15 70007 0 1 400 0 0 z
2 21 15 7000f 1 35 f006 19 20
2 22 16 f000f 1 1 4 0 0 b
2 23 16 b000b 1 1 4 0 0 a
2 24 16 b000f 1 8 20044 22 23 1 0 2
2 25 16 70007 0 1 400 0 0 c
2 26 16 7000f 1 35 f006 24 25
1 a 0 8 7 1 0 2
1 b 0 9 7 1 0 2
1 c 0 10 10008 1 0 2
1 z 0 11 10009 1 0 2
4 21 21 21
4 26 26 26
3 0 adder1 main.add.bit2 ./lib/adder1.v 1 18
2 27 15 f000f 3 1 c 0 0 b
2 28 15 b000b 1 1 4 0 0 a
2 29 15 b000f 3 2 200cc 27 28 1 0 1102
2 30 15 70007 0 1 400 0 0 z
2 31 15 7000f 3 35 f00e 29 30
2 32 16 f000f 3 1 c 0 0 b
2 33 16 b000b 1 1 4 0 0 a
2 34 16 b000f 3 8 200c4 32 33 1 0 2
2 35 16 70007 0 1 400 0 0 c
2 36 16 7000f 1 35 f006 34 35
1 a 0 8 7 1 0 2
1 b 0 9 7 1 0 1102
1 c 0 10 10008 1 0 2
1 z 0 11 10009 1 0 1102
4 31 31 31
4 36 36 36
3 0 adder1 main.add.bit3 ./lib/adder1.v 1 18
2 37 15 f000f 2 1 c 0 0 b
2 38 15 b000b 2 1 c 0 0 a
2 39 15 b000f 3 2 2034c 37 38 1 0 1102
2 40 15 70007 0 1 400 0 0 z
2 41 15 7000f 3 35 f00e 39 40
2 42 16 f000f 2 1 c 0 0 b
2 43 16 b000b 2 1 c 0 0 a
2 44 16 b000f 3 8 2034c 42 43 1 0 102
2 45 16 70007 0 1 400 0 0 c
2 46 16 7000f 2 35 f00e 44 45
1 a 0 8 7 1 0 102
1 b 0 9 7 1 0 102
1 c 0 10 10008 1 0 102
1 z 0 11 10009 1 0 1102
4 41 41 41
4 46 46 46
*/

/* OUTPUT instance2.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : instance2.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    instance2.v                1/    0/    1      100%
  adder4                  adder4.v                   0/    0/    0      100%
  adder1                  adder1.v                   2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    instance2.v                9/    9/   18       50%             8/   10/   18       44%
  adder4                  adder4.v                   6/   10/   16       38%             5/   11/   16       31%
  adder1                  adder1.v                   4/    0/    4      100%             2/    2/    4       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: instance2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h8
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'hc
      ......................... 1->0: 4'h5 ...
      z                         0->1: 4'hc
      ......................... 1->0: 4'hd ...
      carry                     0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      result                    0->1: 5'h1c
      ......................... 1->0: 5'h0d ...

    Module: adder4, File: ./lib/adder4.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h8
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'hc
      ......................... 1->0: 4'h5 ...
      c                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      z                         0->1: 4'hc
      ......................... 1->0: 4'hd ...
      c0                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: adder1, File: ./lib/adder1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              instance2.v                         1/   1/   2       50%
  adder4                            adder4.v                            0/   0/   0      100%
  adder1                            adder1.v                            8/   0/   8      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: instance2.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    assign result = {carry,  z }
                                    |----1-----|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - {}
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    instance2.v               0/   0/   0      100%            0/   0/   0      100%
  adder4                  adder4.v                  0/   0/   0      100%            0/   0/   0      100%
  adder1                  adder1.v                  0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT instance2.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : instance2.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    instance2.v                1/    0/    1      100%
  adder4                  adder4.v                   0/    0/    0      100%
  adder1                  adder1.v                   2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    instance2.v                9/    9/   18       50%             8/   10/   18       44%
  adder4                  adder4.v                   6/   10/   16       38%             5/   11/   16       31%
  adder1                  adder1.v                   4/    0/    4      100%             2/    2/    4       50%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: instance2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h8
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'hc
      ......................... 1->0: 4'h5 ...
      z                         0->1: 4'hc
      ......................... 1->0: 4'hd ...
      carry                     0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      result                    0->1: 5'h1c
      ......................... 1->0: 5'h0d ...

    Module: adder4, File: ./lib/adder4.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h8
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'hc
      ......................... 1->0: 4'h5 ...
      c                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      z                         0->1: 4'hc
      ......................... 1->0: 4'hd ...
      c0                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: adder1, File: ./lib/adder1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              instance2.v                         1/   1/   2       50%
  adder4                            adder4.v                            0/   0/   0      100%
  adder1                            adder1.v                            8/   0/   8      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: instance2.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    assign result = {carry,  z }
                                    |----1-----|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - {}
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    instance2.v               0/   0/   0      100%            0/   0/   0      100%
  adder4                  adder4.v                  0/   0/   0      100%            0/   0/   0      100%
  adder1                  adder1.v                  0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT instance2.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : instance2.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/    0/    1      100%
  <NA>.main.add                                      0/    0/    0      100%
  <NA>.main.add.bit0                                 2/    0/    2      100%
  <NA>.main.add.bit1                                 2/    0/    2      100%
  <NA>.main.add.bit2                                 2/    0/    2      100%
  <NA>.main.add.bit3                                 2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    9/   18       50%             8/   10/   18       44%
  <NA>.main.add                                      6/   10/   16       38%             5/   11/   16       31%
  <NA>.main.add.bit0                                 0/    4/    4        0%             2/    2/    4       50%
  <NA>.main.add.bit1                                 0/    4/    4        0%             0/    4/    4        0%
  <NA>.main.add.bit2                                 2/    2/    4       50%             2/    2/    4       50%
  <NA>.main.add.bit3                                 4/    0/    4      100%             1/    3/    4       25%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: instance2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h8
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'hc
      ......................... 1->0: 4'h5 ...
      z                         0->1: 4'hc
      ......................... 1->0: 4'hd ...
      carry                     0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      result                    0->1: 5'h1c
      ......................... 1->0: 5'h0d ...

    Module: adder4, File: ./lib/adder4.v, Instance: <NA>.main.add
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h8
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'hc
      ......................... 1->0: 4'h5 ...
      c                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      z                         0->1: 4'hc
      ......................... 1->0: 4'hd ...
      c0                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit0
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      z                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit1
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      z                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit2
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit3
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             1/   1/   2       50%
  <NA>.main.add                                                         0/   0/   0      100%
  <NA>.main.add.bit0                                                    4/   4/   8       50%
  <NA>.main.add.bit1                                                    2/   6/   8       25%
  <NA>.main.add.bit2                                                    4/   4/   8       50%
  <NA>.main.add.bit3                                                    6/   2/   8       75%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: instance2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    assign result = {carry,  z }
                                    |----1-----|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - {}
         E | E
        =0=|=1=
         *    


    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit0
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    assign  z  = ( a  ^  b )
                                 |----1----|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    assign  c  = ( a  &  b )
                                 |----1----|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *


    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit1
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    assign  z  = ( a  ^  b )
                                 |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    assign  c  = ( a  &  b )
                                 |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *


    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit2
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    assign  z  = ( a  ^  b )
                                 |----1----|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    assign  c  = ( a  &  b )
                                 |----1----|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *


    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit3
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    assign  z  = ( a  ^  b )
                                 |----1----|

        Expression 1   (3/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *          

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    assign  c  = ( a  &  b )
                                 |----1----|

        Expression 1   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *          



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add                                     0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add.bit0                                0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add.bit1                                0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add.bit2                                0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add.bit3                                0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT instance2.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : instance2.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/    0/    1      100%
  <NA>.main.add                                      0/    0/    0      100%
  <NA>.main.add.bit0                                 2/    0/    2      100%
  <NA>.main.add.bit1                                 2/    0/    2      100%
  <NA>.main.add.bit2                                 2/    0/    2      100%
  <NA>.main.add.bit3                                 2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    9/   18       50%             8/   10/   18       44%
  <NA>.main.add                                      6/   10/   16       38%             5/   11/   16       31%
  <NA>.main.add.bit0                                 0/    4/    4        0%             2/    2/    4       50%
  <NA>.main.add.bit1                                 0/    4/    4        0%             0/    4/    4        0%
  <NA>.main.add.bit2                                 2/    2/    4       50%             2/    2/    4       50%
  <NA>.main.add.bit3                                 4/    0/    4      100%             1/    3/    4       25%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: instance2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h8
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'hc
      ......................... 1->0: 4'h5 ...
      z                         0->1: 4'hc
      ......................... 1->0: 4'hd ...
      carry                     0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      result                    0->1: 5'h1c
      ......................... 1->0: 5'h0d ...

    Module: adder4, File: ./lib/adder4.v, Instance: <NA>.main.add
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h8
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'hc
      ......................... 1->0: 4'h5 ...
      c                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      z                         0->1: 4'hc
      ......................... 1->0: 4'hd ...
      c0                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit0
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      z                         0->1: 1'h0
      ......................... 1->0: 1'h1 ...

    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit1
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      z                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit2
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit3
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             1/   1/   2       50%
  <NA>.main.add                                                         0/   0/   0      100%
  <NA>.main.add.bit0                                                    4/   4/   8       50%
  <NA>.main.add.bit1                                                    2/   6/   8       25%
  <NA>.main.add.bit2                                                    4/   4/   8       50%
  <NA>.main.add.bit3                                                    6/   2/   8       75%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: instance2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    assign result = {carry,  z }
                                    |----1-----|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - {}
         E | E
        =0=|=1=
         *    


    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit0
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    assign  z  = ( a  ^  b )
                                 |----1----|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    assign  c  = ( a  &  b )
                                 |----1----|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *


    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit1
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    assign  z  = ( a  ^  b )
                                 |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    assign  c  = ( a  &  b )
                                 |----1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *


    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit2
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    assign  z  = ( a  ^  b )
                                 |----1----|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    assign  c  = ( a  &  b )
                                 |----1----|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
                   *    *


    Module: adder1, File: ./lib/adder1.v, Instance: <NA>.main.add.bit3
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    assign  z  = ( a  ^  b )
                                 |----1----|

        Expression 1   (3/4)
        ^^^^^^^^^^^^^ - ^
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *          

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    assign  c  = ( a  &  b )
                                 |----1----|

        Expression 1   (3/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *          



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add                                     0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add.bit0                                0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add.bit1                                0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add.bit2                                0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.add.bit3                                0/   0/   0      100%            0/   0/   0      100%


*/
