module main;

parameter STATE_IDLE = 2'b00,
          STATE_HEAD = 2'b01,
          STATE_DATA = 2'b10,
	  STATE_TAIL = 2'b11;

reg            clock;
reg            reset;
reg  [2:0]     state;
reg  [1:0]     next_state;
wire           msg_ip;
reg            head;
reg            tail;
reg            valid;

always @(posedge clock) state <= reset ? {STATE_IDLE,1'b0} : {next_state,(next_state != STATE_IDLE)};

(* covered_fsm, channel, is="state[2:1]", os="next_state" *)
always @(state or head or valid or tail)
  begin
   case( state[2:1] )
     STATE_IDLE:  next_state = (valid & head) ? STATE_HEAD : STATE_IDLE;
     STATE_HEAD:  next_state = (valid & tail) ? STATE_TAIL : STATE_DATA;
     STATE_DATA:  next_state = (valid & tail) ? STATE_TAIL : STATE_DATA;
     STATE_TAIL:  next_state = (valid & head) ? STATE_HEAD : STATE_IDLE;
   endcase
  end

assign msg_ip = state[0];

initial begin
	$dumpfile( "fsm8.1.vcd" );
	$dumpvars( 0, main );
	reset = 1'b1;
	valid = 1'b0;
	head  = 1'b0;
	tail  = 1'b0;
	#20;
	reset = 1'b0;
	@(posedge clock);
        head  <= 1'b1;
        valid <= 1'b1;
	@(posedge clock);
	head  <= 1'b0;
	tail  <= 1'b1;
	@(posedge clock);
	tail  <= 1'b0;
	valid <= 1'b0;
	#20;
	$finish;
end

initial begin
	clock = 1'b0;
	forever #(1) clock = ~clock;
end

endmodule

/* HEADER
GROUPS fsm8.1 all iv vcd lxt
SIM    fsm8.1 all iv vcd  : iverilog fsm8.1.v; ./a.out                             : fsm8.1.vcd
SIM    fsm8.1 all iv lxt  : iverilog fsm8.1.v; ./a.out -lxt2; mv fsm8.1.vcd fsm8.1.lxt : fsm8.1.lxt
SCORE  fsm8.1.vcd     : -t main -vcd fsm8.1.vcd -o fsm8.1.cdd -v fsm8.1.v : fsm8.1.cdd
SCORE  fsm8.1.lxt     : -t main -lxt fsm8.1.lxt -o fsm8.1.cdd -v fsm8.1.v : fsm8.1.cdd
REPORT fsm8.1.cdd 1   : -d v -o fsm8.1.rptM fsm8.1.cdd                         : fsm8.1.rptM
REPORT fsm8.1.cdd 2   : -d v -w -o fsm8.1.rptWM fsm8.1.cdd                     : fsm8.1.rptWM
REPORT fsm8.1.cdd 3   : -d v -i -o fsm8.1.rptI fsm8.1.cdd                      : fsm8.1.rptI
REPORT fsm8.1.cdd 4   : -d v -w -i -o fsm8.1.rptWI fsm8.1.cdd                  : fsm8.1.rptWI
*/

/* OUTPUT fsm8.1.cdd
5 1 * 6 0 0 0 0
3 0 main main fsm8.1.v 1 59
2 1 17 580061 1 32 4 0 0 #STATE_IDLE
2 2 17 4a0053 5 1 c 0 0 next_state
2 3 17 4a0061 6 15 2014c 1 2 1 0 1102
2 4 17 3e0047 5 1 c 0 0 next_state
2 5 17 3e0062 6 31 2024c 3 4 3 0 772a
2 6 17 3d0063 6 26 2000c 5 0 3 0 772a
2 7 17 350038 1 0 20004 0 0 1 1 0
2 8 17 2a0033 1 32 4 0 0 #STATE_IDLE
2 9 17 2a0038 1 31 20044 7 8 33 0 aa aa aa aa aa aa aa aa 2
2 10 17 290039 1 26 20004 9 0 33 0 aa aa aa aa aa aa aa aa 2
2 11 17 210039 7 1a 200cc 6 10 33 0 77aa aa aa aa aa aa aa aa 2
2 12 17 210025 2 1 c 0 0 reset
2 13 17 210063 7 19 201cc 11 12 3 0 772a
2 14 17 18001c 0 1 400 0 0 state
2 15 17 180063 17 38 600e 13 14
2 16 17 110015 2e 1 c 0 0 clock
2 17 17 9000f 0 2a 20000 0 0 2 0 a
2 18 17 90015 46 27 2100a 16 17 1 0 2
2 19 23 3d0046 1 32 4 0 0 #STATE_IDLE
2 20 23 300039 1 32 8 0 0 #STATE_HEAD
2 21 23 1f0039 3 1a 2010c 19 20 32 0 11aa aa aa aa aa aa aa aa
2 22 23 28002b 3 1 c 0 0 head
2 23 23 200024 3 1 c 0 0 valid
2 24 23 20002b 3 8 2024c 22 23 1 0 1102
2 25 23 1f0046 3 19 2024c 21 24 2 0 110a
2 26 23 12001b 0 1 400 0 0 next_state
2 27 23 120046 3 37 600e 25 26
2 28 24 3d0046 1 32 8 0 0 #STATE_DATA
2 29 24 300039 1 32 8 0 0 #STATE_TAIL
2 30 24 1f0039 1 1a 20208 28 29 32 0 aa aa aa aa aa aa aa aa
2 31 24 28002b 1 1 18 0 0 tail
2 32 24 200024 1 1 18 0 0 valid
2 33 24 20002b 1 8 20238 31 32 1 0 2
2 34 24 1f0046 1 19 20238 30 33 2 0 a
2 35 24 12001b 0 1 400 0 0 next_state
2 36 24 120046 1 37 602a 34 35
2 37 25 3d0046 0 32 10 0 0 #STATE_DATA
2 38 25 300039 0 32 10 0 0 #STATE_TAIL
2 39 25 1f0039 0 1a 20030 37 38 32 0 aa aa aa aa aa aa aa aa
2 40 25 28002b 0 1 10 0 0 tail
2 41 25 200024 0 1 10 0 0 valid
2 42 25 20002b 0 8 20030 40 41 1 0 2
2 43 25 1f0046 0 19 20030 39 42 2 0 a
2 44 25 12001b 0 1 400 0 0 next_state
2 45 25 120046 0 37 6022 43 44
2 46 26 3d0046 1 32 4 0 0 #STATE_IDLE
2 47 26 300039 1 32 8 0 0 #STATE_HEAD
2 48 26 1f0039 1 1a 20104 46 47 32 0 aa aa aa aa aa aa aa aa
2 49 26 28002b 1 1 4 0 0 head
2 50 26 200024 1 1 4 0 0 valid
2 51 26 20002b 1 8 20044 49 50 1 0 2
2 52 26 1f0046 1 19 20044 48 51 2 0 a
2 53 26 12001b 0 1 400 0 0 next_state
2 54 26 120046 1 37 6006 52 53
2 55 26 5000e 1 32 8 0 0 #STATE_TAIL
2 56 22 110011 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 57 22 f000f 5 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 58 22 90012 d 24 20e 56 57 state
2 59 26 0 2 2d 2420e 55 58 1 0 102
2 60 25 5000e 1 32 8 0 0 #STATE_DATA
2 61 25 0 2 2d 20206 60 58 1 0 2
2 62 24 5000e 1 32 8 0 0 #STATE_HEAD
2 63 24 0 3 2d 2020e 62 58 1 0 1102
2 64 23 5000e 1 32 4 0 0 #STATE_IDLE
2 65 23 0 6 2d 2014e 64 58 1 0 1102
2 66 20 230026 3 1 c 0 0 tail
2 67 20 230026 0 2a 20000 0 0 2 0 110a
2 68 20 230026 3 29 20008 66 67 1 0 2
2 69 20 1a001e 3 1 c 0 0 valid
2 70 20 1a001e 0 2a 20000 0 0 2 0 110a
2 71 20 1a001e 3 29 20008 69 70 1 0 2
2 72 20 120015 3 1 c 0 0 head
2 73 20 120015 0 2a 20000 0 0 2 0 110a
2 74 20 120015 3 29 20008 72 73 1 0 2
2 75 20 9000d 5 1 c 0 0 state
2 76 20 9000d 0 2a 20000 0 0 4 0 77aa
2 77 20 9000d 5 29 20008 75 76 1 0 2
2 78 20 90015 6 2b 20008 74 77 1 0 2
2 79 20 9001e 6 2b 20008 71 78 1 0 2
2 80 20 90026 d 2b 2100a 68 79 1 0 2
2 81 30 160016 6 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 82 30 100017 6 23 c 0 81 state
2 83 30 7000c 0 1 400 0 0 msg_ip
2 84 30 70017 6 35 f00e 82 83
2 85 55 9000c 1 0 20004 0 0 1 1 0
2 86 55 10005 0 1 400 0 0 clock
2 87 55 1000c 1 37 1006 85 86
2 88 56 17001b 2d 1 1c 0 0 clock
2 89 56 160016 2d 1b 2002c 88 0 1 0 1102
2 90 56 e0012 0 1 400 0 0 clock
2 91 56 e001b 2d 37 602e 89 90
2 92 56 b000b 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 93 56 b000b 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 94 56 9000c 5b 2c 2000a 92 93 32 0 aa aa aa aa aa aa aa aa
2 95 0 0 5 1 f00e 0 0 next_state
2 96 0 0 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 97 0 0 6 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 98 0 0 6 24 f20e 96 97 state
1 #STATE_IDLE 0 0 0 32 0 0 0 0 0 0 0 0 0
1 #STATE_HEAD 0 0 0 32 0 1 0 0 0 0 0 0 0
1 #STATE_DATA 0 0 0 32 0 4 0 0 0 0 0 0 0
1 #STATE_TAIL 0 0 0 32 0 5 0 0 0 0 0 0 0
1 clock 0 8 3000f 1 16 1102
1 reset 0 9 3000f 1 0 1002
1 state 0 10 3000f 3 0 772a
1 next_state 0 11 3000f 2 16 330a
1 msg_ip 0 12 3000f 1 0 1102
1 head 0 13 3000f 1 0 1102
1 tail 0 14 3000f 1 0 1102
1 valid 0 15 3000f 1 0 1102
4 98 98 98
4 95 95 95
4 15 18 18
4 18 15 0
4 54 80 80
4 59 54 80
4 45 80 80
4 61 45 59
4 36 80 80
4 63 36 61
4 27 80 80
4 65 27 63
4 80 65 0
4 84 84 84
4 91 94 94
4 94 91 0
4 87 94 94
6 98 95 1 02,04,04,,01,21,e1,8101
*/

/* OUTPUT fsm8.1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm8.1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm8.1.v                   9/    1/   10       90%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm8.1.v                  10/    1/   11       91%            11/    0/   11      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm8.1.v                           29/  16/  45       64%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm8.1.v                  3/  ? /  ?        ? %            4/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state[2:1]), output state (next_state)

        Hit States

          States
          ======
          2'h0
          2'h1
          2'h3

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      
          2'h0       -> 2'h1      
          2'h1       -> 2'h3      
          2'h3       -> 2'h0      



*/

/* OUTPUT fsm8.1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm8.1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm8.1.v                   9/    1/   10       90%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm8.1.v                  10/    1/   11       91%            11/    0/   11      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm8.1.v                           29/  16/  45       64%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm8.1.v                  3/  ? /  ?        ? %            4/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state[2:1]), output state (next_state)

        Hit States

          States
          ======
          2'h0
          2'h1
          2'h3

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      
          2'h0       -> 2'h1      
          2'h1       -> 2'h3      
          2'h3       -> 2'h0      



*/

/* OUTPUT fsm8.1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm8.1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    1/   10       90%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         10/    1/   11       91%            11/    0/   11      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            29/  16/  45       64%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         3/  ? /  ?        ? %            4/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state[2:1]), output state (next_state)

        Hit States

          States
          ======
          2'h0
          2'h1
          2'h3

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      
          2'h0       -> 2'h1      
          2'h1       -> 2'h3      
          2'h3       -> 2'h0      



*/

/* OUTPUT fsm8.1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm8.1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    1/   10       90%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         10/    1/   11       91%            11/    0/   11      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            29/  16/  45       64%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         3/  ? /  ?        ? %            4/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm8.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state[2:1]), output state (next_state)

        Hit States

          States
          ======
          2'h0
          2'h1
          2'h3

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      
          2'h0       -> 2'h1      
          2'h1       -> 2'h3      
          2'h3       -> 2'h0      



*/
