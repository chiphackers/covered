module main;

reg [const_func(4)-1:0] a;

foo bar[const_func(4)-1:0] (
  .a(a)
);

initial begin
        $dumpfile( "static_func2.vcd" );
        $dumpvars( 0, main );
        #10;
        $finish;
end

function [31:0] const_func;
  input [31:0] size;
  begin
    const_func = 0;
    const_func[size] = 1;
  end
endfunction

endmodule


module foo ( input wire a );

wire b = ~a;

endmodule

/* HEADER
GROUPS static_func2 all vcs vcd
SIM    static_func2 all vcs vcd : vcs +v2k static_func2.v; ./simv                                 : static_func2.vcd
SCORE  static_func2.vcd     : -t main -vcd static_func2.vcd -o static_func2.cdd -v static_func2.v : static_func2.cdd
SCORE  static_func2.lxt     : -t main -lxt static_func2.lxt -o static_func2.cdd -v static_func2.v : static_func2.cdd
REPORT static_func2.cdd 1   : -d v -o static_func2.rptM static_func2.cdd                         : static_func2.rptM
REPORT static_func2.cdd 2   : -d v -w -o static_func2.rptWM static_func2.cdd                     : static_func2.rptWM
REPORT static_func2.cdd 3   : -d v -i -o static_func2.rptI static_func2.cdd                      : static_func2.rptI
REPORT static_func2.cdd 4   : -d v -w -i -o static_func2.rptWI static_func2.cdd                  : static_func2.rptWI
*/

/* OUTPUT static_func2.cdd
5 1 * 6 0 0 0 0
3 0 main main static_func2.v 1 24
1 a 0 3 30018 16 0 aa aa aa aa
3 0 foo main.bar[0] static_func2.v 27 31
2 1 29 a000a 1 1 0 0 0 a
2 2 29 90009 1 1b 20000 1 0 1 0 2
2 3 29 50005 0 1 400 0 0 b
2 4 29 5000a 1 36 f002 2 3
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 4 4 4
3 0 foo main.bar[1] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[2] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[3] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[4] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[5] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[6] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[7] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[8] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[9] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[10] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[11] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[12] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[13] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[14] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 0 foo main.bar[15] static_func2.v 27 31
2 21 29 a000a 1 1 0 0 0 a
2 22 29 90009 1 1b 20000 21 0 1 0 2
2 23 29 50005 0 1 400 0 0 b
2 24 29 5000a 1 36 f002 22 23
1 a 0 27 18 1 0 2
1 b 0 29 30005 1 0 2
4 24 24 24
3 2 main.const_func main.const_func static_func2.v 16 22
2 65 19 110011 0 0 20810 0 0 32 64 0 0 0 0 0 0 0 0
2 66 19 4000d 0 1 c00 0 0 const_func
2 67 19 40011 2 37 11826 65 66
2 68 20 170017 0 0 20810 0 0 32 64 1 0 0 0 0 0 0 0
2 69 20 f0012 0 1 c00 0 0 size
2 70 20 40013 0 23 c00 0 69 const_func
2 71 20 40017 2 37 82a 68 70
1 const_func 0 16 50010 32 16 aa 11aa aa aa aa aa aa aa
1 size 0 17 f 32 16 aa aa aa aa aa aa aa aa
4 71 0 0
4 67 71 71
*/

/* OUTPUT static_func2.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : static_func2.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.v             0/    0/    0      100%
  foo                     static_func2.v             1/    0/    1      100%
  main.const_func         static_func2.v             2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.v             0/   16/   16        0%             0/   16/   16        0%
  foo                     static_func2.v             0/    2/    2        0%             0/    2/    2        0%
  main.const_func         static_func2.v             1/   63/   64        2%             1/   63/   64        2%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 16'h0000
      ......................... 1->0: 16'h0000 ...

    Module: foo, File: static_func2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Function: main.const_func, File: static_func2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      const_func                0->1: 32'h0000_0010
      ......................... 1->0: 32'h0000_0010 ...
      size                      0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              static_func2.v                      0/   0/   0      100%
  foo                               static_func2.v                      0/   2/   2        0%
  main.const_func                   static_func2.v                      0/   0/   0      100%
---------------------------------------------------------------------------------------------------------------------

    Module: foo, File: static_func2.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.v            0/   0/   0      100%            0/   0/   0      100%
  foo                     static_func2.v            0/   0/   0      100%            0/   0/   0      100%
  main.const_func         static_func2.v            0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT static_func2.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : static_func2.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.v             0/    0/    0      100%
  foo                     static_func2.v             1/    0/    1      100%
  main.const_func         static_func2.v             2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.v             0/   16/   16        0%             0/   16/   16        0%
  foo                     static_func2.v             0/    2/    2        0%             0/    2/    2        0%
  main.const_func         static_func2.v             1/   63/   64        2%             1/   63/   64        2%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 16'h0000
      ......................... 1->0: 16'h0000 ...

    Module: foo, File: static_func2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Function: main.const_func, File: static_func2.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      const_func                0->1: 32'h0000_0010
      ......................... 1->0: 32'h0000_0010 ...
      size                      0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              static_func2.v                      0/   0/   0      100%
  foo                               static_func2.v                      0/   2/   2        0%
  main.const_func                   static_func2.v                      0/   0/   0      100%
---------------------------------------------------------------------------------------------------------------------

    Module: foo, File: static_func2.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    static_func2.v            0/   0/   0      100%            0/   0/   0      100%
  foo                     static_func2.v            0/   0/   0      100%            0/   0/   0      100%
  main.const_func         static_func2.v            0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT static_func2.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : static_func2.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%
  <NA>.main.bar[0]                                   1/    0/    1      100%
  <NA>.main.bar[1]                                   1/    0/    1      100%
  <NA>.main.bar[2]                                   1/    0/    1      100%
  <NA>.main.bar[3]                                   1/    0/    1      100%
  <NA>.main.bar[4]                                   1/    0/    1      100%
  <NA>.main.bar[5]                                   1/    0/    1      100%
  <NA>.main.bar[6]                                   1/    0/    1      100%
  <NA>.main.bar[7]                                   1/    0/    1      100%
  <NA>.main.bar[8]                                   1/    0/    1      100%
  <NA>.main.bar[9]                                   1/    0/    1      100%
  <NA>.main.bar[10]                                  1/    0/    1      100%
  <NA>.main.bar[11]                                  1/    0/    1      100%
  <NA>.main.bar[12]                                  1/    0/    1      100%
  <NA>.main.bar[13]                                  1/    0/    1      100%
  <NA>.main.bar[14]                                  1/    0/    1      100%
  <NA>.main.bar[15]                                  1/    0/    1      100%
  <NA>.main.const_func                               2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/   16/   16        0%             0/   16/   16        0%
  <NA>.main.bar[0]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[1]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[2]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[3]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[4]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[5]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[6]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[7]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[8]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[9]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[10]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[11]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[12]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[13]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[14]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[15]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.const_func                               1/   63/   64        2%             1/   63/   64        2%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 16'h0000
      ......................... 1->0: 16'h0000 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[0]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[1]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[2]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[3]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[4]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[5]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[6]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[7]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[8]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[9]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[10]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[11]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[12]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[13]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[14]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[15]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Function: main.const_func, File: static_func2.v, Instance: <NA>.main.const_func
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      const_func                0->1: 32'h0000_0010
      ......................... 1->0: 32'h0000_0010 ...
      size                      0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%
  <NA>.main.bar[0]                                                      0/   2/   2        0%
  <NA>.main.bar[1]                                                      0/   2/   2        0%
  <NA>.main.bar[2]                                                      0/   2/   2        0%
  <NA>.main.bar[3]                                                      0/   2/   2        0%
  <NA>.main.bar[4]                                                      0/   2/   2        0%
  <NA>.main.bar[5]                                                      0/   2/   2        0%
  <NA>.main.bar[6]                                                      0/   2/   2        0%
  <NA>.main.bar[7]                                                      0/   2/   2        0%
  <NA>.main.bar[8]                                                      0/   2/   2        0%
  <NA>.main.bar[9]                                                      0/   2/   2        0%
  <NA>.main.bar[10]                                                     0/   2/   2        0%
  <NA>.main.bar[11]                                                     0/   2/   2        0%
  <NA>.main.bar[12]                                                     0/   2/   2        0%
  <NA>.main.bar[13]                                                     0/   2/   2        0%
  <NA>.main.bar[14]                                                     0/   2/   2        0%
  <NA>.main.bar[15]                                                     0/   2/   2        0%
  <NA>.main.const_func                                                  0/   0/   0      100%
---------------------------------------------------------------------------------------------------------------------

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[0]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[1]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[2]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[3]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[4]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[5]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[6]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[7]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[8]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[9]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[10]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[11]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[12]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[13]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[14]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[15]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[0]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[1]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[2]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[3]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[4]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[5]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[6]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[7]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[8]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[9]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[10]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[11]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[12]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[13]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[14]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[15]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.const_func                              0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT static_func2.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : static_func2.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%
  <NA>.main.bar[0]                                   1/    0/    1      100%
  <NA>.main.bar[1]                                   1/    0/    1      100%
  <NA>.main.bar[2]                                   1/    0/    1      100%
  <NA>.main.bar[3]                                   1/    0/    1      100%
  <NA>.main.bar[4]                                   1/    0/    1      100%
  <NA>.main.bar[5]                                   1/    0/    1      100%
  <NA>.main.bar[6]                                   1/    0/    1      100%
  <NA>.main.bar[7]                                   1/    0/    1      100%
  <NA>.main.bar[8]                                   1/    0/    1      100%
  <NA>.main.bar[9]                                   1/    0/    1      100%
  <NA>.main.bar[10]                                  1/    0/    1      100%
  <NA>.main.bar[11]                                  1/    0/    1      100%
  <NA>.main.bar[12]                                  1/    0/    1      100%
  <NA>.main.bar[13]                                  1/    0/    1      100%
  <NA>.main.bar[14]                                  1/    0/    1      100%
  <NA>.main.bar[15]                                  1/    0/    1      100%
  <NA>.main.const_func                               2/    0/    2      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/   16/   16        0%             0/   16/   16        0%
  <NA>.main.bar[0]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[1]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[2]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[3]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[4]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[5]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[6]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[7]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[8]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[9]                                   0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[10]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[11]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[12]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[13]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[14]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.bar[15]                                  0/    2/    2        0%             0/    2/    2        0%
  <NA>.main.const_func                               1/   63/   64        2%             1/   63/   64        2%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: static_func2.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 16'h0000
      ......................... 1->0: 16'h0000 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[0]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[1]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[2]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[3]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[4]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[5]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[6]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[7]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[8]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[9]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[10]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[11]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[12]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[13]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[14]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[15]
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...

    Function: main.const_func, File: static_func2.v, Instance: <NA>.main.const_func
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      const_func                0->1: 32'h0000_0010
      ......................... 1->0: 32'h0000_0010 ...
      size                      0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%
  <NA>.main.bar[0]                                                      0/   2/   2        0%
  <NA>.main.bar[1]                                                      0/   2/   2        0%
  <NA>.main.bar[2]                                                      0/   2/   2        0%
  <NA>.main.bar[3]                                                      0/   2/   2        0%
  <NA>.main.bar[4]                                                      0/   2/   2        0%
  <NA>.main.bar[5]                                                      0/   2/   2        0%
  <NA>.main.bar[6]                                                      0/   2/   2        0%
  <NA>.main.bar[7]                                                      0/   2/   2        0%
  <NA>.main.bar[8]                                                      0/   2/   2        0%
  <NA>.main.bar[9]                                                      0/   2/   2        0%
  <NA>.main.bar[10]                                                     0/   2/   2        0%
  <NA>.main.bar[11]                                                     0/   2/   2        0%
  <NA>.main.bar[12]                                                     0/   2/   2        0%
  <NA>.main.bar[13]                                                     0/   2/   2        0%
  <NA>.main.bar[14]                                                     0/   2/   2        0%
  <NA>.main.bar[15]                                                     0/   2/   2        0%
  <NA>.main.const_func                                                  0/   0/   0      100%
---------------------------------------------------------------------------------------------------------------------

    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[0]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[1]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[2]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[3]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[4]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[5]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[6]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[7]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[8]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[9]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[10]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[11]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[12]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[13]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[14]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *


    Module: foo, File: static_func2.v, Instance: <NA>.main.bar[15]
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:     b  = ~ a 
                          |1-|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ~
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[0]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[1]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[2]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[3]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[4]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[5]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[6]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[7]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[8]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[9]                                  0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[10]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[11]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[12]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[13]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[14]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.bar[15]                                 0/   0/   0      100%            0/   0/   0      100%
  <NA>.main.const_func                              0/   0/   0      100%            0/   0/   0      100%


*/
