module main;

reg coreclk, sreset, bfr_wr, ld_bfr_data;
reg [31:0] bfr_rd_addr, bfr_wr_addr;

always @(posedge coreclk) begin

  if (sreset)
    bfr_wr_addr <= 3'b0;
  else if (bfr_wr)
    bfr_wr_addr <= bfr_wr_addr + 1'b1;
  else
    bfr_wr_addr <= bfr_wr_addr;

  if (sreset)
    bfr_rd_addr <= 3'b0;
  else if (ld_bfr_data)
    bfr_rd_addr <= bfr_rd_addr + 1'b1;
  else
    bfr_rd_addr <= bfr_rd_addr;

end

initial begin
        $dumpfile( "elseif1.vcd" );
        $dumpvars( 0, main );
	sreset  = 1'b1;
	coreclk = 1'b0;
	#5;
	coreclk = 1'b1;
	#5;
	coreclk = 1'b0;
        #10;
        $finish;
end

endmodule

/* HEADER
GROUPS elseif1 all iv vcs vcd lxt
SIM    elseif1 all iv vcd  : iverilog elseif1.v; ./a.out                             : elseif1.vcd
SIM    elseif1 all iv lxt  : iverilog elseif1.v; ./a.out -lxt2; mv elseif1.vcd elseif1.lxt : elseif1.lxt
SIM    elseif1 all vcs vcd : vcs elseif1.v; ./simv                                   : elseif1.vcd
SCORE  elseif1.vcd     : -t main -vcd elseif1.vcd -o elseif1.cdd -v elseif1.v : elseif1.cdd
SCORE  elseif1.lxt     : -t main -lxt elseif1.lxt -o elseif1.cdd -v elseif1.v : elseif1.cdd
REPORT elseif1.cdd   : -d v -o elseif1.rptM elseif1.cdd                         : elseif1.rptM
REPORT elseif1.cdd   : -d v -w -o elseif1.rptWM elseif1.cdd                     : elseif1.rptWM
REPORT elseif1.cdd   : -d v -i -o elseif1.rptI elseif1.cdd                      : elseif1.rptI
REPORT elseif1.cdd   : -d v -w -i -o elseif1.rptWI elseif1.cdd                  : elseif1.rptWI
*/

/* OUTPUT elseif1.cdd
5 1 * 6 0 0 0 0
3 0 main main elseif1.v 1 37
2 1 9 130016 1 0 20004 0 0 3 1 0
2 2 9 4000e 0 1 400 0 0 bfr_wr_addr
2 3 9 40016 1 38 6006 1 2
2 4 11 210024 0 0 20010 0 0 1 1 1
2 5 11 13001d 0 1 10 0 0 bfr_wr_addr
2 6 11 130024 0 6 20030 4 5 32 0 aa aa aa aa aa aa aa aa
2 7 11 4000e 0 1 400 0 0 bfr_wr_addr
2 8 11 40024 0 38 6022 6 7
2 9 13 13001d 0 1 10 0 0 bfr_wr_addr
2 10 13 4000e 0 1 400 0 0 bfr_wr_addr
2 11 13 4001d 0 38 22 9 10
2 12 10 b0010 0 1 10 0 0 bfr_wr
2 13 10 70011 0 39 22 12 0
2 14 8 6000b 1 1 8 0 0 sreset
2 15 8 2000c 1 39 a 14 0
2 16 16 130016 1 0 20004 0 0 3 1 0
2 17 16 4000e 0 1 400 0 0 bfr_rd_addr
2 18 16 40016 1 38 6006 16 17
2 19 18 210024 0 0 20010 0 0 1 1 1
2 20 18 13001d 0 1 10 0 0 bfr_rd_addr
2 21 18 130024 0 6 20030 19 20 32 0 aa aa aa aa aa aa aa aa
2 22 18 4000e 0 1 400 0 0 bfr_rd_addr
2 23 18 40024 0 38 6022 21 22
2 24 20 13001d 0 1 10 0 0 bfr_rd_addr
2 25 20 4000e 0 1 400 0 0 bfr_rd_addr
2 26 20 4001d 0 38 6022 24 25
2 27 17 b0015 0 1 10 0 0 ld_bfr_data
2 28 17 70016 0 39 22 27 0
2 29 15 6000b 1 1 8 0 0 sreset
2 30 15 2000c 1 39 a 29 0
2 31 6 110017 3 1 c 0 0 coreclk
2 32 6 9000f 0 2a 20000 0 0 2 0 a
2 33 6 90017 5 27 2100a 31 32 1 0 2
1 coreclk 0 3 30004 1 0 1102
1 sreset 0 3 3000d 1 0 2
1 bfr_wr 0 3 30015 1 0 2
1 ld_bfr_data 0 3 3001d 1 0 2
1 bfr_rd_addr 0 4 3000b 32 0 aa aa aa aa aa aa aa aa
1 bfr_wr_addr 0 4 30018 32 0 aa aa aa aa aa aa aa aa
4 26 33 33
4 23 33 33
4 28 23 26
4 18 33 33
4 30 18 28
4 11 30 30
4 8 30 30
4 13 8 11
4 3 30 30
4 15 3 13
4 33 15 0
*/

/* OUTPUT elseif1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : elseif1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    elseif1.v                  5/    6/   11       45%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           10:    if( bfr_wr )
           11:    bfr_wr_addr <= (bfr_wr_addr + 1'b1)
           13:    bfr_wr_addr <= bfr_wr_addr
           17:    if( ld_bfr_data )
           18:    bfr_rd_addr <= (bfr_rd_addr + 1'b1)
           20:    bfr_rd_addr <= bfr_rd_addr



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    elseif1.v                  1/   67/   68        1%             1/   67/   68        1%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      sreset                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bfr_wr                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ld_bfr_data               0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bfr_rd_addr               0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...
      bfr_wr_addr               0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              elseif1.v                           3/  18/  21       14%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              8:    if( sreset )
                        |-1--|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    if( bfr_wr )
                        |-1--|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:    bfr_wr_addr <= (bfr_wr_addr + 1'b1)
                                   |--------1---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             13:    bfr_wr_addr <= bfr_wr_addr
                                   |----1----|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    if( sreset )
                        |-1--|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             17:    if( ld_bfr_data )
                        |----1----|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             18:    bfr_rd_addr <= (bfr_rd_addr + 1'b1)
                                   |--------1---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             20:    bfr_rd_addr <= bfr_rd_addr
                                   |----1----|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    elseif1.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT elseif1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : elseif1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    elseif1.v                  5/    6/   11       45%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           10:    if( bfr_wr )
           11:    bfr_wr_addr <= (bfr_wr_addr + 1'b1)
           13:    bfr_wr_addr <= bfr_wr_addr
           17:    if( ld_bfr_data )
           18:    bfr_rd_addr <= (bfr_rd_addr + 1'b1)
           20:    bfr_rd_addr <= bfr_rd_addr



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    elseif1.v                  1/   67/   68        1%             1/   67/   68        1%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      sreset                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bfr_wr                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ld_bfr_data               0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bfr_rd_addr               0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...
      bfr_wr_addr               0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              elseif1.v                           3/  18/  21       14%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              8:    if( sreset )
                        |-1--|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    if( bfr_wr )
                        |-1--|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:    bfr_wr_addr <= (bfr_wr_addr + 1'b1)
                                   |--------1---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             13:    bfr_wr_addr <= bfr_wr_addr
                                   |----1----|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    if( sreset )
                        |-1--|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             17:    if( ld_bfr_data )
                        |----1----|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             18:    bfr_rd_addr <= (bfr_rd_addr + 1'b1)
                                   |--------1---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             20:    bfr_rd_addr <= bfr_rd_addr
                                   |----1----|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    elseif1.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT elseif1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : elseif1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          5/    6/   11       45%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           10:    if( bfr_wr )
           11:    bfr_wr_addr <= (bfr_wr_addr + 1'b1)
           13:    bfr_wr_addr <= bfr_wr_addr
           17:    if( ld_bfr_data )
           18:    bfr_rd_addr <= (bfr_rd_addr + 1'b1)
           20:    bfr_rd_addr <= bfr_rd_addr



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/   67/   68        1%             1/   67/   68        1%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      sreset                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bfr_wr                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ld_bfr_data               0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bfr_rd_addr               0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...
      bfr_wr_addr               0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             3/  18/  21       14%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              8:    if( sreset )
                        |-1--|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    if( bfr_wr )
                        |-1--|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:    bfr_wr_addr <= (bfr_wr_addr + 1'b1)
                                   |--------1---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             13:    bfr_wr_addr <= bfr_wr_addr
                                   |----1----|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    if( sreset )
                        |-1--|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             17:    if( ld_bfr_data )
                        |----1----|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             18:    bfr_rd_addr <= (bfr_rd_addr + 1'b1)
                                   |--------1---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             20:    bfr_rd_addr <= bfr_rd_addr
                                   |----1----|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT elseif1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : elseif1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          5/    6/   11       45%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           10:    if( bfr_wr )
           11:    bfr_wr_addr <= (bfr_wr_addr + 1'b1)
           13:    bfr_wr_addr <= bfr_wr_addr
           17:    if( ld_bfr_data )
           18:    bfr_rd_addr <= (bfr_rd_addr + 1'b1)
           20:    bfr_rd_addr <= bfr_rd_addr



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/   67/   68        1%             1/   67/   68        1%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      sreset                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bfr_wr                    0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ld_bfr_data               0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bfr_rd_addr               0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...
      bfr_wr_addr               0->1: 32'h0000_0000
      ......................... 1->0: 32'h0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             3/  18/  21       14%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: elseif1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              8:    if( sreset )
                        |-1--|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    if( bfr_wr )
                        |-1--|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:    bfr_wr_addr <= (bfr_wr_addr + 1'b1)
                                   |--------1---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             13:    bfr_wr_addr <= bfr_wr_addr
                                   |----1----|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             15:    if( sreset )
                        |-1--|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             17:    if( ld_bfr_data )
                        |----1----|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             18:    bfr_rd_addr <= (bfr_rd_addr + 1'b1)
                                   |--------1---------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             20:    bfr_rd_addr <= bfr_rd_addr
                                   |----1----|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
