module main;

`define WIDTH  4
`define VALUE  10

wire   [`WIDTH-1:0] a, b, c, d;
reg    [`WIDTH-1:0] e;

assign d = 'd10 + e;
assign c = `WIDTH'd10 + e;
assign b = `WIDTH'd`VALUE + e;
assign a = 'd`VALUE + e;

initial begin
	$dumpfile( "define3.vcd" );
	$dumpvars( 0, main );
	e = `WIDTH'd2;
	#5;
	e = `WIDTH'd3;
	#5;
	$finish;
end

endmodule

/* HEADER
GROUPS define3 all iv vcs vcd lxt
SIM    define3 all iv vcd  : iverilog define3.v; ./a.out                             : define3.vcd
SIM    define3 all iv lxt  : iverilog define3.v; ./a.out -lxt2; mv define3.vcd define3.lxt : define3.lxt
SIM    define3 all vcs vcd : vcs define3.v; ./simv                                   : define3.vcd
SCORE  define3.vcd     : -t main -vcd define3.vcd -o define3.cdd -v define3.v : define3.cdd
SCORE  define3.lxt     : -t main -lxt define3.lxt -o define3.cdd -v define3.v : define3.cdd
REPORT define3.cdd 1   : -d v -o define3.rptM define3.cdd                         : define3.rptM
REPORT define3.cdd 2   : -d v -w -o define3.rptWM define3.cdd                     : define3.rptWM
REPORT define3.cdd 3   : -d v -i -o define3.rptI define3.cdd                      : define3.rptI
REPORT define3.cdd 4   : -d v -w -i -o define3.rptWI define3.cdd                  : define3.rptWI
*/

/* OUTPUT define3.cdd
5 1 * 6 0 0 0 0
3 0 main main define3.v 1 24
2 1 9 120012 2 1 8 0 0 e
2 2 9 b000e 1 0 20008 0 0 32 0 44 0 0 0 0 0 0 0
2 3 9 b0012 3 6 20208 1 2 4 0 1aa
2 4 9 70007 0 1 400 0 0 d
2 5 9 70012 3 35 f00a 3 4
2 6 10 130013 2 1 8 0 0 e
2 7 10 b000f 1 0 20008 0 0 4 0 44
2 8 10 b0013 3 6 20208 6 7 4 0 1aa
2 9 10 70007 0 1 400 0 0 c
2 10 10 70013 3 35 f00a 8 9
2 11 11 130013 2 1 8 0 0 e
2 12 11 b000f 1 0 20008 0 0 4 0 44
2 13 11 b0013 3 6 20208 11 12 4 0 1aa
2 14 11 70007 0 1 400 0 0 b
2 15 11 70013 3 35 f00a 13 14
2 16 12 120012 2 1 8 0 0 e
2 17 12 b000e 1 0 20008 0 0 32 0 44 0 0 0 0 0 0 0
2 18 12 b0012 3 6 20208 16 17 4 0 1aa
2 19 12 70007 0 1 400 0 0 a
2 20 12 70012 3 35 f00a 18 19
1 a 0 6 3000f 4 0 1aa
1 b 0 6 30012 4 0 1aa
1 c 0 6 30015 4 0 1aa
1 d 0 6 30018 4 0 1aa
1 e 0 7 3000f 4 0 1aa
4 5 5 5
4 10 10 10
4 15 15 15
4 20 20 20
*/

/* OUTPUT define3.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : define3.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    define3.v                  4/    0/    4      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    define3.v                  5/   15/   20       25%             0/   20/   20        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: define3.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      c                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      d                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      e                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              define3.v                           4/  12/  16       25%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: define3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    assign  d  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    assign  c  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:    assign  b  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             12:    assign  a  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    define3.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT define3.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : define3.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    define3.v                  4/    0/    4      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    define3.v                  5/   15/   20       25%             0/   20/   20        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: define3.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      c                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      d                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      e                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              define3.v                           4/  12/  16       25%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: define3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    assign  d  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    assign  c  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:    assign  b  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             12:    assign  a  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    define3.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT define3.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : define3.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          4/    0/    4      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          5/   15/   20       25%             0/   20/   20        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: define3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      c                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      d                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      e                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             4/  12/  16       25%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: define3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    assign  d  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    assign  c  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:    assign  b  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             12:    assign  a  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT define3.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : define3.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          4/    0/    4      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          5/   15/   20       25%             0/   20/   20        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: define3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      a                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      b                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      c                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      d                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...
      e                         0->1: 4'h1
      ......................... 1->0: 4'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             4/  12/  16       25%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: define3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
              9:    assign  d  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             10:    assign  c  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             11:    assign  b  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             12:    assign  a  = (10 +  e )
                                 |---1----|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - +
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
