module main;

parameter A       = 0;
parameter STATE_A = 1 << A;

parameter B       = 1;
parameter STATE_B = 1 << B;

parameter C       = 2;
parameter STATE_C = 1 << C;

reg         clock;
reg   [2:0] display_tagto_current_state;
//reg   [2:0] st;
reg   [2:0] next_st;
reg   [7:0] pcix_pio_timeout_recorder;
wire        split_resp_active;
wire  [2:0] split_resp_tag;
reg   [2:0] tag_timeout;
wire        clr_tag_toed;
reg  [79:0] ascii_display_tagto_state;


always @(display_tagto_current_state
//always @(st
   or   pcix_pio_timeout_recorder
   or   split_resp_active
   or   split_resp_tag
   or   tag_timeout
   or   clr_tag_toed) begin // {
    next_st = display_tagto_current_state;
   // next_st = st;
   case(1'b1) // synopsys parallel_case full_case

   //---------------------------------------------------------
   // Idle state: Wait till there is at least one tag timeout.
   //---------------------------------------------------------
   display_tagto_current_state[A]: begin // {
   // st[A]: begin // {
      // synopsys translate_off
      ascii_display_tagto_state = "STATE_A";
      // synopsys translate_on

      if (|pcix_pio_timeout_recorder)
         next_st = STATE_B;
   end // }

   //---------------------------------------------------------
   // Show state: Signal to the rest of the ckty that there is
   // a tag that has timed out. This is a pulse of one pcixclk.
   //---------------------------------------------------------
   display_tagto_current_state[B]: begin // {
   // st[B]: begin // {
      // synopsys translate_off
      ascii_display_tagto_state = "STATE_B";
      // synopsys translate_on

      next_st = STATE_C;
   end // }

   //---------------------------------------------------------
   // No Show state: Wait until all the reuired actions have
   // been taken for the tag that has timed out.
   //---------------------------------------------------------
   display_tagto_current_state[C]: begin // {
   // st[C]: begin // {
      // synopsys translate_off
      ascii_display_tagto_state = "STATE_C";
      // synopsys translate_on

      if (clr_tag_toed
      ||  (split_resp_active && (split_resp_tag == tag_timeout)))
         next_st = STATE_A;
   end // }
   endcase
end // }

always @(posedge clock) display_tagto_current_state <= next_st;
// always @(posedge clock) st <= next_st;

initial begin
	$dumpfile( "case4.1.vcd" );
	$dumpvars( 0, main );
	#50;
	$finish;
end

initial begin
	clock = 1'b0;
	forever #(1) clock = ~clock;
end

endmodule

/* HEADER
GROUPS case4.1 all iv vcs vcd lxt
SIM    case4.1 all iv vcd  : iverilog case4.1.v; ./a.out                             : case4.1.vcd
SIM    case4.1 all iv lxt  : iverilog case4.1.v; ./a.out -lxt2; mv case4.1.vcd case4.1.lxt : case4.1.lxt
SIM    case4.1 all vcs vcd : vcs case4.1.v; ./simv                                   : case4.1.vcd
SCORE  case4.1.vcd     : -t main -vcd case4.1.vcd -o case4.1.cdd -v case4.1.v : case4.1.cdd
SCORE  case4.1.lxt     : -t main -lxt case4.1.lxt -o case4.1.cdd -v case4.1.v : case4.1.cdd
REPORT case4.1.cdd 1   : -d v -o case4.1.rptM case4.1.cdd                         : case4.1.rptM
REPORT case4.1.cdd 2   : -d v -w -o case4.1.rptWM case4.1.cdd                     : case4.1.rptWM
REPORT case4.1.cdd 3   : -d v -i -o case4.1.rptI case4.1.cdd                      : case4.1.rptI
REPORT case4.1.cdd 4   : -d v -w -i -o case4.1.rptWI case4.1.cdd                  : case4.1.rptWI
*/

/* OUTPUT case4.1.cdd
5 1 * 6 0 0 0 0
3 0 main main case4.1.v 1 93
2 1 31 e0028 1 1 0 0 0 display_tagto_current_state
2 2 31 4000a 0 1 400 0 0 next_st
2 3 31 40028 1 37 2 1 2
2 4 41 22002a 0 0 20010 0 0 56 4 1 10 55 11 11 10 10 11 1 10 10 11 5 11
2 5 41 6001e 0 1 400 0 0 ascii_display_tagto_state
2 6 41 6002a 0 37 22 4 5
2 7 45 130019 0 32 10 0 0 #STATE_B
2 8 45 9000f 0 1 400 0 0 next_st
2 9 45 90019 0 37 6022 7 8
2 10 44 b0023 0 1 10 0 0 pcix_pio_timeout_recorder
2 11 44 a000a 0 1e 20020 10 0 1 0 2
2 12 44 60024 0 39 4022 11 0
2 13 55 22002a 0 0 20010 0 0 56 4 4 10 55 11 11 10 10 11 1 10 10 11 5 11
2 14 55 6001e 0 1 400 0 0 ascii_display_tagto_state
2 15 55 6002a 0 37 22 13 14
2 16 58 100016 0 32 10 0 0 #STATE_C
2 17 58 6000c 0 1 400 0 0 next_st
2 18 58 60016 0 37 6022 16 17
2 19 68 22002a 0 0 20010 0 0 56 4 5 10 55 11 11 10 10 11 1 10 10 11 5 11
2 20 68 6001e 0 1 400 0 0 ascii_display_tagto_state
2 21 68 6002a 0 37 22 19 20
2 22 73 130019 0 32 10 0 0 #STATE_A
2 23 73 9000f 0 1 400 0 0 next_st
2 24 73 90019 0 37 6022 22 23
2 25 72 33003d 0 1 10 0 0 tag_timeout
2 26 72 21002e 0 1 10 0 0 split_resp_tag
2 27 72 21003d 0 11 20030 25 26 1 0 2
2 28 72 b001b 0 1 10 0 0 split_resp_active
2 29 72 b003e 0 18 20030 27 28 1 0 2
2 30 71 a0015 0 1 10 0 0 clr_tag_toed
2 31 71 a003f 0 17 20030 29 30 1 0 2
2 32 71 60040 0 39 4022 31 0
2 33 65 1f001f 1 32 8 0 0 #C
2 34 65 30020 1 23 0 0 33 display_tagto_current_state
2 35 33 8000b 3 0 2000a 0 0 1 1 1
2 36 65 0 1 2d 24006 34 35 1 0 2
2 37 52 1f001f 1 32 8 0 0 #B
2 38 52 30020 1 23 0 0 37 display_tagto_current_state
2 39 52 0 1 2d 20006 38 35 1 0 2
2 40 38 1f001f 1 32 4 0 0 #A
2 41 38 30020 1 23 0 0 40 display_tagto_current_state
2 42 38 0 1 2d 20006 41 35 1 0 2
2 43 30 80013 1 1 0 0 0 clr_tag_toed
2 44 30 80013 0 2a 20000 0 0 2 0 a
2 45 30 80013 1 29 20008 43 44 1 0 2
2 46 29 80012 1 1 0 0 0 tag_timeout
2 47 29 80012 0 2a 20000 0 0 4 0 aa
2 48 29 80012 1 29 20000 46 47 1 0 2
2 49 28 80015 1 1 0 0 0 split_resp_tag
2 50 28 80015 0 2a 20000 0 0 4 0 aa
2 51 28 80015 1 29 20008 49 50 1 0 2
2 52 27 80018 1 1 0 0 0 split_resp_active
2 53 27 80018 0 2a 20000 0 0 2 0 a
2 54 27 80018 1 29 20008 52 53 1 0 2
2 55 26 80020 1 1 0 0 0 pcix_pio_timeout_recorder
2 56 26 80020 0 2a 20000 0 0 9 0 aa aa 2
2 57 26 80020 1 29 20000 55 56 1 0 2
2 58 24 90023 1 1 0 0 0 display_tagto_current_state
2 59 24 90023 0 2a 20000 0 0 4 0 aa
2 60 24 90023 1 29 20000 58 59 1 0 2
2 61 24 90020 1 2b 20000 57 60 1 0 2
2 62 24 90018 1 2b 20008 54 61 1 0 2
2 63 24 90015 1 2b 20008 51 62 1 0 2
2 64 24 90012 1 2b 20008 48 63 1 0 2
2 65 24 90013 3 2b 2100a 45 64 1 0 2
2 66 78 37003d 1 1 0 0 0 next_st
2 67 78 180032 0 1 400 0 0 display_tagto_current_state
2 68 78 18003d 19 38 6002 66 67
2 69 78 110015 33 1 c 0 0 clock
2 70 78 9000f 0 2a 20000 0 0 2 0 a
2 71 78 90015 4d 27 2100a 69 70 1 0 2
2 72 89 9000c 1 0 20004 0 0 1 1 0
2 73 89 10005 0 1 400 0 0 clock
2 74 89 1000c 1 37 1006 72 73
2 75 90 17001b 32 1 1c 0 0 clock
2 76 90 160016 32 1b 2002c 75 0 1 0 1102
2 77 90 e0012 0 1 400 0 0 clock
2 78 90 e001b 32 37 602e 76 77
2 79 90 b000b 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 80 90 b000b 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 81 90 9000c 65 2c 2000a 79 80 32 0 aa aa aa aa aa aa aa aa
1 #A 0 0 0 32 0 0 0 0 0 0 0 0 0
1 #STATE_A 0 0 0 32 0 101 0 0 0 0 0 0 0
1 #B 0 0 0 32 0 1 0 0 0 0 0 0 0
1 #STATE_B 0 0 0 32 0 204 0 0 0 0 0 0 0
1 #C 0 0 0 32 0 4 0 0 0 0 0 0 0
1 #STATE_C 0 0 0 32 0 410 0 0 0 0 0 0 0
1 clock 0 12 3000c 1 16 1102
1 display_tagto_current_state 0 13 3000c 3 0 2a
1 next_st 0 15 3000c 3 16 2a
1 pcix_pio_timeout_recorder 0 16 3000c 8 0 aa aa
1 split_resp_active 0 17 3000c 1 0 2
1 split_resp_tag 0 18 3000c 3 0 2a
1 tag_timeout 0 19 3000c 3 0 2a
1 clr_tag_toed 0 20 3000c 1 0 2
1 ascii_display_tagto_state 0 21 3000c 80 16 aa aa aa aa aa aa aa aa aa aa aa aa aa aa aa aa aa aa aa aa
4 24 65 65
4 32 24 65
4 21 32 32
4 36 21 65
4 18 65 65
4 15 18 18
4 39 15 36
4 9 65 65
4 12 9 65
4 6 12 12
4 42 6 39
4 3 42 42
4 65 3 0
4 68 71 71
4 71 68 0
4 78 81 81
4 81 78 0
4 74 81 81
*/

/* OUTPUT case4.1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : case4.1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.1.v                  6/    8/   14       43%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           41:    ascii_display_tagto_state = "STATE_A"
           44:    if( |pcix_pio_timeout_recorder )
           45:    next_st = STATE_B
           55:    ascii_display_tagto_state = "STATE_B"
           58:    next_st = STATE_C
           68:    ascii_display_tagto_state = "STATE_C"
           71:    if( (clr_tag_toed || ...
           73:    next_st = STATE_A



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.1.v                  1/  102/  103        1%             1/  102/  103        1%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      display_tagto_current_state  0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      next_st                   0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      pcix_pio_timeout_recorder  0->1: 8'h00
      ......................... 1->0: 8'h00 ...
      split_resp_active         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      split_resp_tag            0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      tag_timeout               0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      clr_tag_toed              0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ascii_display_tagto_state  0->1: 80'h0000_0000_0000_0000_0000
      ......................... 1->0: 80'h0000_0000_0000_0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              case4.1.v                           6/  19/  25       24%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    @(display_tagto_current_state or 
                      |------------1------------|    
                    pcix_pio_timeout_recorder or 
                    |-----------2-----------|    
                    split_resp_active or 
                    split_resp_tag or 
                    tag_timeout or 
                    |----3----|    
                    clr_tag_toed)

        Expression 1   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

        Expression 2   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

        Expression 3   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    next_st = display_tagto_current_state
                              |------------1------------|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             44:    if( |pcix_pio_timeout_recorder )
                        |-----------1------------|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - |
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             71:    if( (clr_tag_toed || 
                        |-------3---------
                    (split_resp_active && (split_resp_tag == tag_timeout))) )
                                          |--------------1--------------|    
                    |-------------------------2--------------------------|   
                    ---------------------------3--------------------------|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 2   (0/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 3   (0/4)
        ^^^^^^^^^^^^^ - ||
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    display_tagto_current_state <= next_st
                                                   |--1--|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.1.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT case4.1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : case4.1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.1.v                  6/    8/   14       43%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           41:    ascii_display_tagto_state = "STATE_A"
           44:    if( |pcix_pio_timeout_recorder )
           45:    next_st = STATE_B
           55:    ascii_display_tagto_state = "STATE_B"
           58:    next_st = STATE_C
           68:    ascii_display_tagto_state = "STATE_C"
           71:    if( (clr_tag_toed || (split_resp_active && (split_resp_tag == tag_timeout))) )
           73:    next_st = STATE_A



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.1.v                  1/  102/  103        1%             1/  102/  103        1%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      display_tagto_current_state  0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      next_st                   0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      pcix_pio_timeout_recorder  0->1: 8'h00
      ......................... 1->0: 8'h00 ...
      split_resp_active         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      split_resp_tag            0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      tag_timeout               0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      clr_tag_toed              0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ascii_display_tagto_state  0->1: 80'h0000_0000_0000_0000_0000
      ......................... 1->0: 80'h0000_0000_0000_0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              case4.1.v                           6/  19/  25       24%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    @(display_tagto_current_state or pcix_pio_timeout_recorder or split_resp_active or split_resp_tag or 
                      |------------1------------|    |-----------2-----------|                                           
                    tag_timeout or clr_tag_toed)
                    |----3----|                 

        Expression 1   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

        Expression 2   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

        Expression 3   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    next_st = display_tagto_current_state
                              |------------1------------|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             44:    if( |pcix_pio_timeout_recorder )
                        |-----------1------------|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - |
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             71:    if( (clr_tag_toed || (split_resp_active && (split_resp_tag == tag_timeout))) )
                                                               |--------------1--------------|    
                                         |-------------------------2--------------------------|   
                        |----------------------------------3-----------------------------------|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 2   (0/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 3   (0/4)
        ^^^^^^^^^^^^^ - ||
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    display_tagto_current_state <= next_st
                                                   |--1--|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    case4.1.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT case4.1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : case4.1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          6/    8/   14       43%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           41:    ascii_display_tagto_state = "STATE_A"
           44:    if( |pcix_pio_timeout_recorder )
           45:    next_st = STATE_B
           55:    ascii_display_tagto_state = "STATE_B"
           58:    next_st = STATE_C
           68:    ascii_display_tagto_state = "STATE_C"
           71:    if( (clr_tag_toed || ...
           73:    next_st = STATE_A



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/  102/  103        1%             1/  102/  103        1%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      display_tagto_current_state  0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      next_st                   0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      pcix_pio_timeout_recorder  0->1: 8'h00
      ......................... 1->0: 8'h00 ...
      split_resp_active         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      split_resp_tag            0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      tag_timeout               0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      clr_tag_toed              0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ascii_display_tagto_state  0->1: 80'h0000_0000_0000_0000_0000
      ......................... 1->0: 80'h0000_0000_0000_0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             6/  19/  25       24%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    @(display_tagto_current_state or 
                      |------------1------------|    
                    pcix_pio_timeout_recorder or 
                    |-----------2-----------|    
                    split_resp_active or 
                    split_resp_tag or 
                    tag_timeout or 
                    |----3----|    
                    clr_tag_toed)

        Expression 1   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

        Expression 2   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

        Expression 3   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    next_st = display_tagto_current_state
                              |------------1------------|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             44:    if( |pcix_pio_timeout_recorder )
                        |-----------1------------|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - |
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             71:    if( (clr_tag_toed || 
                        |-------3---------
                    (split_resp_active && (split_resp_tag == tag_timeout))) )
                                          |--------------1--------------|    
                    |-------------------------2--------------------------|   
                    ---------------------------3--------------------------|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 2   (0/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 3   (0/4)
        ^^^^^^^^^^^^^ - ||
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    display_tagto_current_state <= next_st
                                                   |--1--|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT case4.1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : case4.1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          6/    8/   14       43%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           41:    ascii_display_tagto_state = "STATE_A"
           44:    if( |pcix_pio_timeout_recorder )
           45:    next_st = STATE_B
           55:    ascii_display_tagto_state = "STATE_B"
           58:    next_st = STATE_C
           68:    ascii_display_tagto_state = "STATE_C"
           71:    if( (clr_tag_toed || (split_resp_active && (split_resp_tag == tag_timeout))) )
           73:    next_st = STATE_A



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          1/  102/  103        1%             1/  102/  103        1%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      display_tagto_current_state  0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      next_st                   0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      pcix_pio_timeout_recorder  0->1: 8'h00
      ......................... 1->0: 8'h00 ...
      split_resp_active         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      split_resp_tag            0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      tag_timeout               0->1: 3'h0
      ......................... 1->0: 3'h0 ...
      clr_tag_toed              0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ascii_display_tagto_state  0->1: 80'h0000_0000_0000_0000_0000
      ......................... 1->0: 80'h0000_0000_0000_0000_0000 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             6/  19/  25       24%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: case4.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    @(display_tagto_current_state or pcix_pio_timeout_recorder or split_resp_active or split_resp_tag or 
                      |------------1------------|    |-----------2-----------|                                           
                    tag_timeout or clr_tag_toed)
                    |----3----|                 

        Expression 1   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

        Expression 2   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

        Expression 3   (0/1)
        ^^^^^^^^^^^^^ - 
         * Event did not occur

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    next_st = display_tagto_current_state
                              |------------1------------|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             44:    if( |pcix_pio_timeout_recorder )
                        |-----------1------------|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - |
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             71:    if( (clr_tag_toed || (split_resp_active && (split_resp_tag == tag_timeout))) )
                                                               |--------------1--------------|    
                                         |-------------------------2--------------------------|   
                        |----------------------------------3-----------------------------------|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *   *

        Expression 2   (0/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 3   (0/4)
        ^^^^^^^^^^^^^ - ||
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             78:    display_tagto_current_state <= next_st
                                                   |--1--|

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
