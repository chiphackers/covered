module main;

reg        clock;
reg        reset;
reg        a, b;
reg [21:0] c, d;

reg [3:0] addr;
reg       wr;

always @(posedge clock)
  begin
   if( reset )
     begin
      a <= 1'b0;
      b <= 1'b0;
      c <= 22'h0;
     end
   else if( (addr == 4'h0) && wr)
     a <= 1'b1;
   else if( (addr == 4'h1) && wr)
     b <= 1'b1;
   else 
     begin
      if( d[ 0] ) c[0]  <= 1'b1;
      if( d[ 1] ) c[1]  <= 1'b1;
      if( d[ 2] ) c[2]  <= 1'b1;
      if( d[ 3] ) c[3]  <= 1'b1;
      if( d[ 4] ) c[4]  <= 1'b1;
      if( d[ 5] ) c[5]  <= 1'b1;
      if( d[ 6] ) c[6]  <= 1'b1;
      if( d[ 7] ) c[7]  <= 1'b1;
      if( d[ 8] ) c[8]  <= 1'b1;
      if( d[ 9] ) c[9]  <= 1'b1;
      if( d[10] ) c[10] <= 1'b1;
      if( d[11] ) c[11] <= 1'b1;
      if( d[12] ) c[12] <= 1'b1;
      if( d[13] ) c[13] <= 1'b1;
      if( d[14] ) c[14] <= 1'b1;
      if( d[15] ) c[15] <= 1'b1;
      if( d[16] ) c[16] <= 1'b1;
      if( d[17] ) c[17] <= 1'b1;
      if( d[18] ) c[18] <= 1'b1;
      if( d[19] ) c[19] <= 1'b1;
      if( d[20] ) c[20] <= 1'b1;
      if( d[21] ) c[21] <= 1'b1;
     end
  end

initial begin
	$dumpfile( "always9.vcd" );
	$dumpvars( 0, main );
	reset = 1'b1;
	addr  = 4'h0;
	d[8]  = 1'b1;
        wr    = 1'b0;
	#20;
	reset = 1'b0;
	#20;
	wr    = 1'b1;
	#20;
	$finish;
end

initial begin
	clock = 1'b0;
	forever #(1) clock = ~clock;
end

endmodule

/* HEADER
GROUPS always9 all iv vcs vcd lxt
SIM    always9 all iv vcd  : iverilog always9.v; ./a.out                             : always9.vcd
SIM    always9 all iv lxt  : iverilog always9.v; ./a.out -lxt2; mv always9.vcd always9.lxt : always9.lxt
SIM    always9 all vcs vcd : vcs always9.v; ./simv                                   : always9.vcd
SCORE  always9.vcd     : -t main -vcd always9.vcd -o always9.cdd -v always9.v : always9.cdd
SCORE  always9.lxt     : -t main -lxt always9.lxt -o always9.cdd -v always9.v : always9.cdd
REPORT always9.cdd 1   : -d v -o always9.rptM always9.cdd                         : always9.rptM
REPORT always9.cdd 2   : -d v -w -o always9.rptWM always9.cdd                     : always9.rptWM
REPORT always9.cdd 3   : -d v -i -o always9.rptI always9.cdd                      : always9.rptI
REPORT always9.cdd 4   : -d v -w -i -o always9.rptWI always9.cdd                  : always9.rptWI
*/

/* OUTPUT always9.cdd
5 1 * 6 0 0 0 0
3 0 main main always9.v 1 70
2 1 15 b000e 1 0 20004 0 0 1 1 0
2 2 15 60006 0 1 400 0 0 a
2 3 15 6000e a 38 6 1 2
2 4 16 b000e 1 0 20004 0 0 1 1 0
2 5 16 60006 0 1 400 0 0 b
2 6 16 6000e a 38 6 4 5
2 7 17 b000f 1 0 20004 0 0 22 3 0 0 0 0 0 0
2 8 17 60006 0 1 400 0 0 c
2 9 17 6000f a 38 6006 7 8
2 10 20 a000d 1 0 20008 0 0 1 1 1
2 11 20 50005 0 1 400 0 0 a
2 12 20 5000d a 38 600a 10 11
2 13 22 a000d 0 0 20010 0 0 1 1 1
2 14 22 50005 0 1 400 0 0 b
2 15 22 5000d 0 38 6022 13 14
2 16 25 1b001e 0 0 20010 0 0 1 1 1
2 17 25 140014 0 0 20400 0 0 32 64 0 0 0 0 0 0 0 0
2 18 25 120015 0 23 400 0 17 c
2 19 25 12001e 0 38 22 16 18
2 20 25 d000d 1 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 21 25 a000e 1 23 0 0 20 d
2 22 25 60010 a 39 4002 21 0
2 23 26 1b001e 0 0 20010 0 0 1 1 1
2 24 26 140014 0 0 20400 0 0 32 64 1 0 0 0 0 0 0 0
2 25 26 120015 0 23 400 0 24 c
2 26 26 12001e 0 38 22 23 25
2 27 26 d000d 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 28 26 a000e 1 23 0 0 27 d
2 29 26 60010 a 39 4002 28 0
2 30 27 1b001e 0 0 20010 0 0 1 1 1
2 31 27 140014 0 0 20400 0 0 32 64 4 0 0 0 0 0 0 0
2 32 27 120015 0 23 400 0 31 c
2 33 27 12001e 0 38 22 30 32
2 34 27 d000d 1 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 35 27 a000e 1 23 0 0 34 d
2 36 27 60010 a 39 4002 35 0
2 37 28 1b001e 0 0 20010 0 0 1 1 1
2 38 28 140014 0 0 20400 0 0 32 64 5 0 0 0 0 0 0 0
2 39 28 120015 0 23 400 0 38 c
2 40 28 12001e 0 38 22 37 39
2 41 28 d000d 1 0 20008 0 0 32 64 5 0 0 0 0 0 0 0
2 42 28 a000e 1 23 0 0 41 d
2 43 28 60010 a 39 4002 42 0
2 44 29 1b001e 0 0 20010 0 0 1 1 1
2 45 29 140014 0 0 20400 0 0 32 64 10 0 0 0 0 0 0 0
2 46 29 120015 0 23 400 0 45 c
2 47 29 12001e 0 38 22 44 46
2 48 29 d000d 1 0 20008 0 0 32 64 10 0 0 0 0 0 0 0
2 49 29 a000e 1 23 0 0 48 d
2 50 29 60010 a 39 4002 49 0
2 51 30 1b001e 0 0 20010 0 0 1 1 1
2 52 30 140014 0 0 20400 0 0 32 64 11 0 0 0 0 0 0 0
2 53 30 120015 0 23 400 0 52 c
2 54 30 12001e 0 38 22 51 53
2 55 30 d000d 1 0 20008 0 0 32 64 11 0 0 0 0 0 0 0
2 56 30 a000e 1 23 0 0 55 d
2 57 30 60010 a 39 4002 56 0
2 58 31 1b001e 0 0 20010 0 0 1 1 1
2 59 31 140014 0 0 20400 0 0 32 64 14 0 0 0 0 0 0 0
2 60 31 120015 0 23 400 0 59 c
2 61 31 12001e 0 38 22 58 60
2 62 31 d000d 1 0 20008 0 0 32 64 14 0 0 0 0 0 0 0
2 63 31 a000e 1 23 0 0 62 d
2 64 31 60010 a 39 4002 63 0
2 65 32 1b001e 0 0 20010 0 0 1 1 1
2 66 32 140014 0 0 20400 0 0 32 64 15 0 0 0 0 0 0 0
2 67 32 120015 0 23 400 0 66 c
2 68 32 12001e 0 38 22 65 67
2 69 32 d000d 1 0 20008 0 0 32 64 15 0 0 0 0 0 0 0
2 70 32 a000e 1 23 0 0 69 d
2 71 32 60010 a 39 4002 70 0
2 72 33 1b001e 1 0 20008 0 0 1 1 1
2 73 33 140014 0 0 20400 0 0 32 64 40 0 0 0 0 0 0 0
2 74 33 120015 0 23 400 0 73 c
2 75 33 12001e a 38 a 72 74
2 76 33 d000d 1 0 20008 0 0 32 64 40 0 0 0 0 0 0 0
2 77 33 a000e 1 23 8 0 76 d
2 78 33 60010 a 39 400a 77 0
2 79 34 1b001e 0 0 20010 0 0 1 1 1
2 80 34 140014 0 0 20400 0 0 32 64 41 0 0 0 0 0 0 0
2 81 34 120015 0 23 400 0 80 c
2 82 34 12001e 0 38 22 79 81
2 83 34 d000d 1 0 20008 0 0 32 64 41 0 0 0 0 0 0 0
2 84 34 a000e 1 23 0 0 83 d
2 85 34 60010 a 39 4002 84 0
2 86 35 1b001e 0 0 20010 0 0 1 1 1
2 87 35 140015 0 0 20400 0 0 32 64 44 0 0 0 0 0 0 0
2 88 35 120016 0 23 400 0 87 c
2 89 35 12001e 0 38 22 86 88
2 90 35 c000d 1 0 20008 0 0 32 64 44 0 0 0 0 0 0 0
2 91 35 a000e 1 23 0 0 90 d
2 92 35 60010 a 39 4002 91 0
2 93 36 1b001e 0 0 20010 0 0 1 1 1
2 94 36 140015 0 0 20400 0 0 32 64 45 0 0 0 0 0 0 0
2 95 36 120016 0 23 400 0 94 c
2 96 36 12001e 0 38 22 93 95
2 97 36 c000d 1 0 20008 0 0 32 64 45 0 0 0 0 0 0 0
2 98 36 a000e 1 23 0 0 97 d
2 99 36 60010 a 39 4002 98 0
2 100 37 1b001e 0 0 20010 0 0 1 1 1
2 101 37 140015 0 0 20400 0 0 32 64 50 0 0 0 0 0 0 0
2 102 37 120016 0 23 400 0 101 c
2 103 37 12001e 0 38 22 100 102
2 104 37 c000d 1 0 20008 0 0 32 64 50 0 0 0 0 0 0 0
2 105 37 a000e 1 23 0 0 104 d
2 106 37 60010 a 39 4002 105 0
2 107 38 1b001e 0 0 20010 0 0 1 1 1
2 108 38 140015 0 0 20400 0 0 32 64 51 0 0 0 0 0 0 0
2 109 38 120016 0 23 400 0 108 c
2 110 38 12001e 0 38 22 107 109
2 111 38 c000d 1 0 20008 0 0 32 64 51 0 0 0 0 0 0 0
2 112 38 a000e 1 23 0 0 111 d
2 113 38 60010 a 39 4002 112 0
2 114 39 1b001e 0 0 20010 0 0 1 1 1
2 115 39 140015 0 0 20400 0 0 32 64 54 0 0 0 0 0 0 0
2 116 39 120016 0 23 400 0 115 c
2 117 39 12001e 0 38 22 114 116
2 118 39 c000d 1 0 20008 0 0 32 64 54 0 0 0 0 0 0 0
2 119 39 a000e 1 23 0 0 118 d
2 120 39 60010 a 39 4002 119 0
2 121 40 1b001e 0 0 20010 0 0 1 1 1
2 122 40 140015 0 0 20400 0 0 32 64 55 0 0 0 0 0 0 0
2 123 40 120016 0 23 400 0 122 c
2 124 40 12001e 0 38 22 121 123
2 125 40 c000d 1 0 20008 0 0 32 64 55 0 0 0 0 0 0 0
2 126 40 a000e 1 23 0 0 125 d
2 127 40 60010 a 39 4002 126 0
2 128 41 1b001e 0 0 20010 0 0 1 1 1
2 129 41 140015 0 0 20400 0 0 32 64 0 1 0 0 0 0 0 0
2 130 41 120016 0 23 400 0 129 c
2 131 41 12001e 0 38 22 128 130
2 132 41 c000d 1 0 20008 0 0 32 64 0 1 0 0 0 0 0 0
2 133 41 a000e 1 23 0 0 132 d
2 134 41 60010 a 39 4002 133 0
2 135 42 1b001e 0 0 20010 0 0 1 1 1
2 136 42 140015 0 0 20400 0 0 32 64 1 1 0 0 0 0 0 0
2 137 42 120016 0 23 400 0 136 c
2 138 42 12001e 0 38 22 135 137
2 139 42 c000d 1 0 20008 0 0 32 64 1 1 0 0 0 0 0 0
2 140 42 a000e 1 23 0 0 139 d
2 141 42 60010 a 39 4002 140 0
2 142 43 1b001e 0 0 20010 0 0 1 1 1
2 143 43 140015 0 0 20400 0 0 32 64 4 1 0 0 0 0 0 0
2 144 43 120016 0 23 400 0 143 c
2 145 43 12001e 0 38 22 142 144
2 146 43 c000d 1 0 20008 0 0 32 64 4 1 0 0 0 0 0 0
2 147 43 a000e 1 23 0 0 146 d
2 148 43 60010 a 39 4002 147 0
2 149 44 1b001e 0 0 20010 0 0 1 1 1
2 150 44 140015 0 0 20400 0 0 32 64 5 1 0 0 0 0 0 0
2 151 44 120016 0 23 400 0 150 c
2 152 44 12001e 0 38 22 149 151
2 153 44 c000d 1 0 20008 0 0 32 64 5 1 0 0 0 0 0 0
2 154 44 a000e 1 23 0 0 153 d
2 155 44 60010 a 39 4002 154 0
2 156 45 1b001e 0 0 20010 0 0 1 1 1
2 157 45 140015 0 0 20400 0 0 32 64 10 1 0 0 0 0 0 0
2 158 45 120016 0 23 400 0 157 c
2 159 45 12001e 0 38 22 156 158
2 160 45 c000d 1 0 20008 0 0 32 64 10 1 0 0 0 0 0 0
2 161 45 a000e 1 23 0 0 160 d
2 162 45 60010 a 39 4002 161 0
2 163 46 1b001e 0 0 20010 0 0 1 1 1
2 164 46 140015 0 0 20400 0 0 32 64 11 1 0 0 0 0 0 0
2 165 46 120016 0 23 400 0 164 c
2 166 46 12001e 0 38 6022 163 165
2 167 46 c000d 1 0 20008 0 0 32 64 11 1 0 0 0 0 0 0
2 168 46 a000e 1 23 0 0 167 d
2 169 46 60010 a 39 4002 168 0
2 170 21 1e001f 1 1 14 0 0 wr
2 171 21 150018 1 0 20008 0 0 4 3 1
2 172 21 d0010 1 1 4 0 0 addr
2 173 21 d0018 1 11 20084 171 172 1 0 2
2 174 21 c001f 1 18 20064 170 173 1 0 2
2 175 21 80020 a 39 26 174 0
2 176 19 1e001f 2 1 c 0 0 wr
2 177 19 150018 1 0 20004 0 0 4 3 0
2 178 19 d0010 1 1 4 0 0 addr
2 179 19 d0018 1 11 20048 177 178 1 0 2
2 180 19 c001f 2 18 2030c 176 179 1 0 102
2 181 19 80020 14 39 e 180 0
2 182 13 7000b 2 1 c 0 0 reset
2 183 13 3000d 1e 39 e 182 0
2 184 11 110015 3d 1 c 0 0 clock
2 185 11 9000f 0 2a 20000 0 0 2 0 a
2 186 11 90015 5c 27 2100a 184 185 1 0 2
2 187 66 9000c 1 0 20004 0 0 1 1 0
2 188 66 10005 0 1 400 0 0 clock
2 189 66 1000c 1 37 1006 187 188
2 190 67 17001b 3c 1 1c 0 0 clock
2 191 67 160016 3c 1b 2002c 190 0 1 0 1102
2 192 67 e0012 0 1 400 0 0 clock
2 193 67 e001b 3c 37 602e 191 192
2 194 67 b000b 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 195 67 b000b 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 196 67 9000c 79 2c 2000a 194 195 32 0 aa aa aa aa aa aa aa aa
1 clock 0 3 3000b 1 16 1102
1 reset 0 4 3000b 1 0 1002
1 a 0 5 3000b 1 0 102
1 b 0 5 3000e 1 0 2
1 c 0 6 3000b 22 0 aa aa 1aa aa aa a
1 d 0 6 3000e 22 0 aa aa aa aa aa a
1 addr 0 8 3000a 4 0 aa
1 wr 0 9 3000a 1 0 102
4 166 186 186
4 169 166 186
4 159 169 169
4 162 159 169
4 152 162 162
4 155 152 162
4 145 155 155
4 148 145 155
4 138 148 148
4 141 138 148
4 131 141 141
4 134 131 141
4 124 134 134
4 127 124 134
4 117 127 127
4 120 117 127
4 110 120 120
4 113 110 120
4 103 113 113
4 106 103 113
4 96 106 106
4 99 96 106
4 89 99 99
4 92 89 99
4 82 92 92
4 85 82 92
4 75 85 85
4 78 75 85
4 68 78 78
4 71 68 78
4 61 71 71
4 64 61 71
4 54 64 64
4 57 54 64
4 47 57 57
4 50 47 57
4 40 50 50
4 43 40 50
4 33 43 43
4 36 33 43
4 26 36 36
4 29 26 36
4 19 29 29
4 22 19 29
4 15 186 186
4 175 15 22
4 12 186 186
4 181 12 175
4 9 186 186
4 6 9 9
4 3 6 6
4 183 3 181
4 186 183 0
4 193 196 196
4 196 193 0
4 189 196 196
*/

/* OUTPUT always9.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : always9.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    always9.v                 33/   22/   55       60%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           22:     b  <= 1'b1
           25:    c[0] <= 1'b1
           26:    c[1] <= 1'b1
           27:    c[2] <= 1'b1
           28:    c[3] <= 1'b1
           29:    c[4] <= 1'b1
           30:    c[5] <= 1'b1
           31:    c[6] <= 1'b1
           32:    c[7] <= 1'b1
           34:    c[9] <= 1'b1
           35:    c[10] <= 1'b1
           36:    c[11] <= 1'b1
           37:    c[12] <= 1'b1
           38:    c[13] <= 1'b1
           39:    c[14] <= 1'b1
           40:    c[15] <= 1'b1
           41:    c[16] <= 1'b1
           42:    c[17] <= 1'b1
           43:    c[18] <= 1'b1
           44:    c[19] <= 1'b1
           45:    c[20] <= 1'b1
           46:    c[21] <= 1'b1



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    always9.v                  4/   49/   53        8%             2/   51/   53        4%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 22'h00_0100
      ......................... 1->0: 22'h00_0000 ...
      d                         0->1: 22'h00_0000
      ......................... 1->0: 22'h00_0000 ...
      addr                      0->1: 4'h0
      ......................... 1->0: 4'h0 ...
      wr                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              always9.v                          11/  50/  61       18%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             19:    if( ((addr == 4'h0) &&  wr) )
                         |-----1------|          
                        |----------2----------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 2   (2/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    if( ((addr == 4'h1) &&  wr) )
                         |-----1------|          
                        |----------2----------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
             *

        Expression 2   (1/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    if( d[0] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    if( d[1] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    if( d[2] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    if( d[3] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    if( d[4] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             30:    if( d[5] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    if( d[6] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             32:    if( d[7] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             33:    if( d[8] )
                        |1-|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             34:    if( d[9] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             35:    if( d[10] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             36:    if( d[11] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             37:    if( d[12] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             38:    if( d[13] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             39:    if( d[14] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             40:    if( d[15] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             41:    if( d[16] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             42:    if( d[17] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             43:    if( d[18] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             44:    if( d[19] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             45:    if( d[20] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             46:    if( d[21] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    always9.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT always9.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : always9.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    always9.v                 33/   22/   55       60%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           22:     b  <= 1'b1
           25:    c[0] <= 1'b1
           26:    c[1] <= 1'b1
           27:    c[2] <= 1'b1
           28:    c[3] <= 1'b1
           29:    c[4] <= 1'b1
           30:    c[5] <= 1'b1
           31:    c[6] <= 1'b1
           32:    c[7] <= 1'b1
           34:    c[9] <= 1'b1
           35:    c[10] <= 1'b1
           36:    c[11] <= 1'b1
           37:    c[12] <= 1'b1
           38:    c[13] <= 1'b1
           39:    c[14] <= 1'b1
           40:    c[15] <= 1'b1
           41:    c[16] <= 1'b1
           42:    c[17] <= 1'b1
           43:    c[18] <= 1'b1
           44:    c[19] <= 1'b1
           45:    c[20] <= 1'b1
           46:    c[21] <= 1'b1



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    always9.v                  4/   49/   53        8%             2/   51/   53        4%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 22'h00_0100
      ......................... 1->0: 22'h00_0000 ...
      d                         0->1: 22'h00_0000
      ......................... 1->0: 22'h00_0000 ...
      addr                      0->1: 4'h0
      ......................... 1->0: 4'h0 ...
      wr                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              always9.v                          11/  50/  61       18%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             19:    if( ((addr == 4'h0) &&  wr) )
                         |-----1------|          
                        |----------2----------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 2   (2/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    if( ((addr == 4'h1) &&  wr) )
                         |-----1------|          
                        |----------2----------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
             *

        Expression 2   (1/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    if( d[0] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    if( d[1] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    if( d[2] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    if( d[3] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    if( d[4] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             30:    if( d[5] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    if( d[6] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             32:    if( d[7] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             33:    if( d[8] )
                        |1-|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             34:    if( d[9] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             35:    if( d[10] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             36:    if( d[11] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             37:    if( d[12] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             38:    if( d[13] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             39:    if( d[14] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             40:    if( d[15] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             41:    if( d[16] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             42:    if( d[17] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             43:    if( d[18] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             44:    if( d[19] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             45:    if( d[20] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             46:    if( d[21] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    always9.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT always9.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : always9.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         33/   22/   55       60%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           22:     b  <= 1'b1
           25:    c[0] <= 1'b1
           26:    c[1] <= 1'b1
           27:    c[2] <= 1'b1
           28:    c[3] <= 1'b1
           29:    c[4] <= 1'b1
           30:    c[5] <= 1'b1
           31:    c[6] <= 1'b1
           32:    c[7] <= 1'b1
           34:    c[9] <= 1'b1
           35:    c[10] <= 1'b1
           36:    c[11] <= 1'b1
           37:    c[12] <= 1'b1
           38:    c[13] <= 1'b1
           39:    c[14] <= 1'b1
           40:    c[15] <= 1'b1
           41:    c[16] <= 1'b1
           42:    c[17] <= 1'b1
           43:    c[18] <= 1'b1
           44:    c[19] <= 1'b1
           45:    c[20] <= 1'b1
           46:    c[21] <= 1'b1



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          4/   49/   53        8%             2/   51/   53        4%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 22'h00_0100
      ......................... 1->0: 22'h00_0000 ...
      d                         0->1: 22'h00_0000
      ......................... 1->0: 22'h00_0000 ...
      addr                      0->1: 4'h0
      ......................... 1->0: 4'h0 ...
      wr                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            11/  50/  61       18%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             19:    if( ((addr == 4'h0) &&  wr) )
                         |-----1------|          
                        |----------2----------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 2   (2/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    if( ((addr == 4'h1) &&  wr) )
                         |-----1------|          
                        |----------2----------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
             *

        Expression 2   (1/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    if( d[0] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    if( d[1] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    if( d[2] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    if( d[3] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    if( d[4] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             30:    if( d[5] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    if( d[6] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             32:    if( d[7] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             33:    if( d[8] )
                        |1-|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             34:    if( d[9] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             35:    if( d[10] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             36:    if( d[11] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             37:    if( d[12] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             38:    if( d[13] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             39:    if( d[14] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             40:    if( d[15] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             41:    if( d[16] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             42:    if( d[17] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             43:    if( d[18] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             44:    if( d[19] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             45:    if( d[20] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             46:    if( d[21] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT always9.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : always9.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         33/   22/   55       60%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           22:     b  <= 1'b1
           25:    c[0] <= 1'b1
           26:    c[1] <= 1'b1
           27:    c[2] <= 1'b1
           28:    c[3] <= 1'b1
           29:    c[4] <= 1'b1
           30:    c[5] <= 1'b1
           31:    c[6] <= 1'b1
           32:    c[7] <= 1'b1
           34:    c[9] <= 1'b1
           35:    c[10] <= 1'b1
           36:    c[11] <= 1'b1
           37:    c[12] <= 1'b1
           38:    c[13] <= 1'b1
           39:    c[14] <= 1'b1
           40:    c[15] <= 1'b1
           41:    c[16] <= 1'b1
           42:    c[17] <= 1'b1
           43:    c[18] <= 1'b1
           44:    c[19] <= 1'b1
           45:    c[20] <= 1'b1
           46:    c[21] <= 1'b1



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          4/   49/   53        8%             2/   51/   53        4%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      a                         0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b                         0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c                         0->1: 22'h00_0100
      ......................... 1->0: 22'h00_0000 ...
      d                         0->1: 22'h00_0000
      ......................... 1->0: 22'h00_0000 ...
      addr                      0->1: 4'h0
      ......................... 1->0: 4'h0 ...
      wr                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            11/  50/  61       18%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: always9.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             19:    if( ((addr == 4'h0) &&  wr) )
                         |-----1------|          
                        |----------2----------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
         *    

        Expression 2   (2/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    if( ((addr == 4'h1) &&  wr) )
                         |-----1------|          
                        |----------2----------|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ==
         E | E
        =0=|=1=
             *

        Expression 2   (1/4)
        ^^^^^^^^^^^^^ - &&
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    if( d[0] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             26:    if( d[1] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             27:    if( d[2] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             28:    if( d[3] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             29:    if( d[4] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             30:    if( d[5] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             31:    if( d[6] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             32:    if( d[7] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             33:    if( d[8] )
                        |1-|  

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             34:    if( d[9] )
                        |1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             35:    if( d[10] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             36:    if( d[11] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             37:    if( d[12] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             38:    if( d[13] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             39:    if( d[14] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             40:    if( d[15] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             41:    if( d[16] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             42:    if( d[17] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             43:    if( d[18] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             44:    if( d[19] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             45:    if( d[20] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             46:    if( d[21] )
                        |-1-|  

        Expression 1   (0/2)
        ^^^^^^^^^^^^^ - []
         E | E
        =0=|=1=
         *   *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
