module main;

integer a;

initial a <<= 2;

endmodule
