module main;

integer a;

initial a--;

endmodule
