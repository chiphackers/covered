module main;

foo f();

endmodule

//---------------------------------

module foo (
  output wire [1:0] a
);

endmodule
