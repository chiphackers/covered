/*
 Name:        null_stmt1.8.v
 Author:      Trevor Williams  (phase1geo@gmail.com)
 Date:        03/13/2008
 Purpose:     Verify that null statements after case statements work properly.
 Simulators:  IV CVER VERIWELL VCS
 Modes:       VCD LXT VPI
*/

module main;

reg a, b;

initial begin
	a = 1'b0;
	b = 1'b0;
	#5;
	case( a )
          1'b0 : ;
          1'b1 : b = 1'b1;
        endcase
	a = 1'b1;
end

initial begin
`ifdef DUMP
        $dumpfile( "null_stmt1.8.vcd" );
        $dumpvars( 0, main );
`endif
        #10;
        $finish;
end

endmodule
