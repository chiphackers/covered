module main;

wire    qo, ro, so, to, uo, vo, wo, xo;

wire    q1, r1, s1, t1, u1, v1;

reg     s2;
reg     t2;
reg     u2;
reg     v2;

reg     w1, w2, w3;
reg     x1, x2, x3;


tran( qo, q1 );
rtran( ro, r1 );
tranif0( so, s1, s2 );
tranif1( to, t1, t2 );
rtranif0( uo, u1, u2 );
rtranif1( vo, v1, v2 );

cmos( wo, w1, w2, w3 );
rcmos( xo, x1, x2, x3 );

initial begin
	$dumpfile( "gate1.1.vcd" );
	$dumpvars( 0, main );
	s2 = 1'b0;
	t2 = 1'b0;
	u2 = 1'b0;
	v2 = 1'b0;
	w1 = 1'b0;
	w2 = 1'b0;
	w3 = 1'b0;
	x1 = 1'b0;
	x2 = 1'b0;
	x3 = 1'b0;
	#5;
	s2 = 1'b1;
	t2 = 1'b1;
	u2 = 1'b1;
	v2 = 1'b1;
	w2 = 1'b1;
	x2 = 1'b1;
	#5;
	$finish;
end

endmodule

/* HEADER
GROUPS gate1.1 all vcs vcd
SIM    gate1.1 all vcs vcd : vcs gate1.1.v; ./simv                                   : gate1.1.vcd
SCORE  gate1.1.vcd     : -t main -vcd gate1.1.vcd -o gate1.1.cdd -v gate1.1.v : gate1.1.cdd
SCORE  gate1.1.lxt     : -t main -lxt gate1.1.lxt -o gate1.1.cdd -v gate1.1.v : gate1.1.cdd
REPORT gate1.1.cdd 1   : -d v -o gate1.1.rptM gate1.1.cdd                         : gate1.1.rptM
REPORT gate1.1.cdd 2   : -d v -w -o gate1.1.rptWM gate1.1.cdd                     : gate1.1.rptWM
REPORT gate1.1.cdd 3   : -d v -i -o gate1.1.rptI gate1.1.cdd                      : gate1.1.rptI
REPORT gate1.1.cdd 4   : -d v -w -i -o gate1.1.rptWI gate1.1.cdd                  : gate1.1.rptWI
*/

/* OUTPUT gate1.1.cdd
5 1 * 6 0 0 0 0
3 0 main main gate1.1.v 1 50
1 qo 0 3 30008 1 0 2
1 ro 0 3 3000c 1 0 2
1 so 0 3 30010 1 0 2
1 to 0 3 30014 1 0 2
1 uo 0 3 30018 1 0 2
1 vo 0 3 3001c 1 0 2
1 wo 0 3 30020 1 0 2
1 xo 0 3 30024 1 0 2
1 q1 0 5 30008 1 0 2
1 r1 0 5 3000c 1 0 2
1 s1 0 5 30010 1 0 2
1 t1 0 5 30014 1 0 2
1 u1 0 5 30018 1 0 2
1 v1 0 5 3001c 1 0 2
1 s2 0 7 30008 1 0 102
1 t2 0 8 30008 1 0 102
1 u2 0 9 30008 1 0 102
1 v2 0 10 30008 1 0 102
1 w1 0 12 30008 1 0 2
1 w2 0 12 3000c 1 0 102
1 w3 0 12 30010 1 0 2
1 x1 0 13 30008 1 0 2
1 x2 0 13 3000c 1 0 102
1 x3 0 13 30010 1 0 2
*/

/* OUTPUT gate1.1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : gate1.1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.1.v                  0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.1.v                  6/   18/   24       25%             0/   24/   24        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: gate1.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      qo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ro                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      so                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      to                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      uo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      vo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      wo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      xo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      q1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      r1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      s1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      t1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      u1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      v1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      s2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      t2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      u2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      v2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      w1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      w2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      w3                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      x3                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              gate1.1.v                           0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.1.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT gate1.1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : gate1.1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.1.v                  0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.1.v                  6/   18/   24       25%             0/   24/   24        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: gate1.1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      qo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ro                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      so                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      to                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      uo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      vo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      wo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      xo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      q1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      r1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      s1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      t1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      u1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      v1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      s2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      t2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      u2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      v2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      w1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      w2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      w3                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      x3                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              gate1.1.v                           0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.1.v                 0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT gate1.1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : gate1.1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          6/   18/   24       25%             0/   24/   24        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: gate1.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      qo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ro                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      so                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      to                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      uo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      vo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      wo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      xo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      q1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      r1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      s1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      t1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      u1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      v1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      s2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      t2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      u2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      v2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      w1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      w2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      w3                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      x3                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT gate1.1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : gate1.1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          6/   18/   24       25%             0/   24/   24        0%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: gate1.1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      qo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ro                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      so                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      to                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      uo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      vo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      wo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      xo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      q1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      r1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      s1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      t1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      u1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      v1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      s2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      t2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      u2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      v2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      w1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      w2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      w3                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x1                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      x2                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      x3                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
