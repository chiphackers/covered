module main;

reg a;

(* foo, bar, pan *)
initial a = 1'b0;

endmodule
