module level3a(
  input  wire a,
  output wire b
);

assign b = a ? 0 : 1;

endmodule
