module main;

wire    ao, bo, co, do, eo, fo, go, ho, io, jo, ko, lo, mo, no, oo, po;

reg     a1, a2;
reg     b1, b2;
reg     c1, c2;
reg     d1, d2;
reg     e1, e2;
reg     f1, f2;

reg     g1;
reg     h1;

reg     i1, i2;
reg     j1, j2;
reg     k1, k2;
reg     l1, l2;

reg     m1, m2;
reg     n1, n2;
reg     o1, o2;
reg     p1, p2;


and( ao, a1, a2 );
nand( bo, b1, b2 );
or( co, c1, c2 );
nor( do, d1, d2 );
xor( eo, e1, e2 );
xnor( fo, f1, f2 );

buf( go, g1 );
not( ho, h1 );

bufif0( io, i1, i2 );
bufif1( jo, j1, j2 );
notif0( ko, k1, k2 );
notif1( lo, l1, l2 );

nmos( mo, m1, m2 );
pmos( no, n1, n2 );
rnmos( oo, o1, o2 );
rpmos( po, p1, p2 );


initial begin
	$dumpfile( "gate1.vcd" );
	$dumpvars( 0, main );
	a1 = 1'b0;
	a2 = 1'b0;
	b1 = 1'b0;
	b2 = 1'b0;
	c1 = 1'b0;
	c2 = 1'b0;
	d1 = 1'b0;
	d2 = 1'b0;
	e1 = 1'b0;
	e2 = 1'b0;
	f1 = 1'b0;
	f2 = 1'b0;
	g1 = 1'b0;
	h1 = 1'b0;
	i1 = 1'b0;
	i2 = 1'b0;
	j1 = 1'b0;
	j2 = 1'b0;
	k1 = 1'b0;
	k2 = 1'b0;
	l1 = 1'b0;
	l2 = 1'b0;
	m1 = 1'b0;
	m2 = 1'b0;
	n1 = 1'b0;
	n2 = 1'b0;
	o1 = 1'b0;
	o2 = 1'b0;
	p1 = 1'b0;
	p2 = 1'b0;
	#5;
	a1 = 1'b1;
	b1 = 1'b1;
	c1 = 1'b1;
	d1 = 1'b1;
	e1 = 1'b1;
	f1 = 1'b1;
	g1 = 1'b1;
	h1 = 1'b1;
	i1 = 1'b1;
	j1 = 1'b1;
	k1 = 1'b1;
	l1 = 1'b1;
	m1 = 1'b1;
	n1 = 1'b1;
	o1 = 1'b1;
	p1 = 1'b1;
	#5;
	$finish;
end

endmodule

/* HEADER
GROUPS gate1 all iv vcs vcd lxt
SIM    gate1 all iv vcd  : iverilog gate1.v; ./a.out                             : gate1.vcd
SIM    gate1 all iv lxt  : iverilog gate1.v; ./a.out -lxt2; mv gate1.vcd gate1.lxt : gate1.lxt
SIM    gate1 all vcs vcd : vcs gate1.v; ./simv                                   : gate1.vcd
SCORE  gate1.vcd     : -t main -vcd gate1.vcd -o gate1.cdd -v gate1.v : gate1.cdd
SCORE  gate1.lxt     : -t main -lxt gate1.lxt -o gate1.cdd -v gate1.v : gate1.cdd
REPORT gate1.cdd 1   : -d v -o gate1.rptM gate1.cdd                         : gate1.rptM
REPORT gate1.cdd 2   : -d v -w -o gate1.rptWM gate1.cdd                     : gate1.rptWM
REPORT gate1.cdd 3   : -d v -i -o gate1.rptI gate1.cdd                      : gate1.rptI
REPORT gate1.cdd 4   : -d v -w -i -o gate1.rptWI gate1.cdd                  : gate1.rptWI
*/

/* OUTPUT gate1.cdd
5 1 * 6 0 0 0 0
3 0 main main gate1.v 1 101
1 ao 0 3 30008 1 0 2
1 bo 0 3 3000c 1 0 2
1 co 0 3 30010 1 0 102
1 do 0 3 30014 1 0 1002
1 eo 0 3 30018 1 0 102
1 fo 0 3 3001c 1 0 1002
1 go 0 3 30020 1 0 102
1 ho 0 3 30024 1 0 1002
1 io 0 3 30028 1 0 102
1 jo 0 3 3002c 1 0 2
1 ko 0 3 30030 1 0 1002
1 lo 0 3 30034 1 0 2
1 mo 0 3 30038 1 0 2
1 no 0 3 3003c 1 0 102
1 oo 0 3 30040 1 0 2
1 po 0 3 30044 1 0 102
1 a1 0 5 30008 1 0 102
1 a2 0 5 3000c 1 0 2
1 b1 0 6 30008 1 0 102
1 b2 0 6 3000c 1 0 2
1 c1 0 7 30008 1 0 102
1 c2 0 7 3000c 1 0 2
1 d1 0 8 30008 1 0 102
1 d2 0 8 3000c 1 0 2
1 e1 0 9 30008 1 0 102
1 e2 0 9 3000c 1 0 2
1 f1 0 10 30008 1 0 102
1 f2 0 10 3000c 1 0 2
1 g1 0 12 30008 1 0 102
1 h1 0 13 30008 1 0 102
1 i1 0 15 30008 1 0 102
1 i2 0 15 3000c 1 0 2
1 j1 0 16 30008 1 0 102
1 j2 0 16 3000c 1 0 2
1 k1 0 17 30008 1 0 102
1 k2 0 17 3000c 1 0 2
1 l1 0 18 30008 1 0 102
1 l2 0 18 3000c 1 0 2
1 m1 0 20 30008 1 0 102
1 m2 0 20 3000c 1 0 2
1 n1 0 21 30008 1 0 102
1 n2 0 21 3000c 1 0 2
1 o1 0 22 30008 1 0 102
1 o2 0 22 3000c 1 0 2
1 p1 0 23 30008 1 0 102
1 p2 0 23 3000c 1 0 2
*/

/* OUTPUT gate1.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : gate1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.v                    0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.v                   22/   24/   46       48%             4/   42/   46        9%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: gate1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      ao                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      co                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      do                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      eo                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      fo                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      ho                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      io                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      jo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ko                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      lo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      mo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      no                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      oo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      po                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      a1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      a2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      d2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      e1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      e2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      f2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      g1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      h1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      i1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      i2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      j1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      j2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      k1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      k2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      l1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      l2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      m1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      m2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      n1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      n2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      o1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      o2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      p1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      p2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              gate1.v                             0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.v                   0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT gate1.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : gate1.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.v                    0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.v                   22/   24/   46       48%             4/   42/   46        9%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: gate1.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      ao                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      co                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      do                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      eo                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      fo                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      ho                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      io                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      jo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ko                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      lo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      mo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      no                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      oo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      po                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      a1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      a2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      d2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      e1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      e2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      f2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      g1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      h1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      i1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      i2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      j1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      j2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      k1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      k2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      l1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      l2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      m1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      m2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      n1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      n2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      o1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      o2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      p1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      p2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              gate1.v                             0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    gate1.v                   0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT gate1.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : gate1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         22/   24/   46       48%             4/   42/   46        9%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: gate1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      ao                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      co                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      do                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      eo                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      fo                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      ho                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      io                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      jo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ko                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      lo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      mo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      no                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      oo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      po                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      a1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      a2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      d2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      e1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      e2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      f2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      g1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      h1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      i1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      i2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      j1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      j2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      k1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      k2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      l1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      l2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      m1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      m2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      n1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      n2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      o1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      o2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      p1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      p2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/

/* OUTPUT gate1.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : gate1.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          0/    0/    0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         22/   24/   46       48%             4/   42/   46        9%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: gate1.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      ao                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      bo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      co                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      do                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      eo                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      fo                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      go                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      ho                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      io                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      jo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      ko                        0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      lo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      mo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      no                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      oo                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      po                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      a1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      a2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      b1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      b2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      c1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      c2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      d1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      d2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      e1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      e2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      f1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      f2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      g1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      h1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      i1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      i2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      j1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      j2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      k1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      k2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      l1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      l2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      m1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      m2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      n1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      n2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      o1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      o2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...
      p1                        0->1: 1'h1
      ......................... 1->0: 1'h0 ...
      p2                        0->1: 1'h0
      ......................... 1->0: 1'h0 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                             0/   0/   0      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         0/   0/   0      100%            0/   0/   0      100%


*/
