module main;

parameter STATE_IDLE = 16'h0001,
          STATE_HEAD = 16'h0010,
          STATE_DATA = 16'h0100,
          STATE_TAIL = 16'h1000;

reg         clk;
reg         reset;
reg         head;
reg         tail;
reg         valid;
reg [15:0]  state;
reg [15:0]  next_state;

always @(posedge clk) state <= reset ? STATE_IDLE : next_state;

always @(state or head or valid or tail)
  begin
   case( state )
     STATE_IDLE:  next_state = (valid & head) ? STATE_HEAD : STATE_IDLE;
     STATE_HEAD:  next_state = (valid & tail) ? STATE_TAIL : STATE_DATA;
     STATE_DATA:  next_state = (valid & tail) ? STATE_TAIL : STATE_DATA;
     STATE_TAIL:  next_state = (valid & head) ? STATE_HEAD : STATE_IDLE;
   endcase
  end

initial begin
	$dumpfile( "fsm3.vcd" );
	$dumpvars( 0, main );
        reset = 1'b1;
	head  = 1'b0;
        tail  = 1'b0;
        valid = 1'b0;
	#20;
	reset = 1'b0;
	#20;
	@(posedge clk);
        head <= 1'b1;
	valid <= 1'b1;
	@(posedge clk);
        head <= 1'b0;
	#20;
	@(posedge clk);
        tail <= 1'b1;
	@(posedge clk);
	tail <= 1'b0;
	head <= 1'b1;
	@(posedge clk);
	tail <= 1'b1;
        head <= 1'b0;
	@(posedge clk);
	tail  <= 1'b0;
	valid <= 1'b0;
	#20;
	$finish;
end

initial begin
	clk = 1'b0;
        forever #(2) clk = ~clk;
end

endmodule

/* HEADER
GROUPS fsm3 all iv vcs vcd lxt
SIM    fsm3 all iv vcd  : iverilog fsm3.v; ./a.out                             : fsm3.vcd
SIM    fsm3 all iv lxt  : iverilog fsm3.v; ./a.out -lxt2; mv fsm3.vcd fsm3.lxt : fsm3.lxt
SIM    fsm3 all vcs vcd : vcs fsm3.v; ./simv                                   : fsm3.vcd
SCORE  fsm3.vcd     : -t main -vcd fsm3.vcd -o fsm3.cdd -y lib -v fsm3.v -F main=state,next_state : fsm3.cdd
SCORE  fsm3.lxt     : -t main -lxt fsm3.lxt -o fsm3.cdd -y lib -v fsm3.v -F main=state,next_state : fsm3.cdd
REPORT fsm3.cdd 1   : -d v -o fsm3.rptM fsm3.cdd                         : fsm3.rptM
REPORT fsm3.cdd 2   : -d v -w -o fsm3.rptWM fsm3.cdd                     : fsm3.rptWM
REPORT fsm3.cdd 3   : -d v -i -o fsm3.rptI fsm3.cdd                      : fsm3.rptI
REPORT fsm3.cdd 4   : -d v -w -i -o fsm3.rptWI fsm3.cdd                  : fsm3.rptWI
*/

/* OUTPUT fsm3.cdd
5 1 * 6 0 0 0 0
3 0 main main fsm3.v 1 64
2 1 16 34003d 9 1 8 0 0 next_state
2 2 16 270030 1 32 8 0 0 #STATE_IDLE
2 3 16 1f0030 b 1a 20208 1 2 32 0 11aa 11aa 11aa 11aa aa aa aa aa
2 4 16 1f0023 2 1 c 0 0 reset
2 5 16 1f003d b 19 20288 3 4 16 0 11aa 11aa 11aa 11aa
2 6 16 16001a 0 1 400 0 0 state
2 7 16 16003d 19 38 600a 5 6
2 8 16 110013 32 1 c 0 0 clk
2 9 16 9000f 0 2a 20000 0 0 2 0 a
2 10 16 90013 4c 27 2100a 8 9 1 0 2
2 11 21 3d0046 1 32 8 0 0 #STATE_IDLE
2 12 21 300039 1 32 8 0 0 #STATE_HEAD
2 13 21 1f0039 3 1a 20208 11 12 32 0 11aa 11aa aa aa aa aa aa aa
2 14 21 28002b 3 1 c 0 0 head
2 15 21 200024 3 1 c 0 0 valid
2 16 21 20002b 3 8 2024c 14 15 1 0 1102
2 17 21 1f0046 3 19 20288 13 16 16 0 11aa 11aa aa aa
2 18 21 12001b 0 1 400 0 0 next_state
2 19 21 120046 3 37 600a 17 18
2 20 22 3d0046 1 32 8 0 0 #STATE_DATA
2 21 22 300039 1 32 8 0 0 #STATE_TAIL
2 22 22 1f0039 2 1a 20208 20 21 32 0 aa aa 10aa 1aa aa aa aa aa
2 23 22 28002b 2 1 1c 0 0 tail
2 24 22 200024 1 1 18 0 0 valid
2 25 22 20002b 2 8 2033c 23 24 1 0 102
2 26 22 1f0046 2 19 202b8 22 25 16 0 aa aa 10aa 1aa
2 27 22 12001b 0 1 400 0 0 next_state
2 28 22 120046 2 37 602a 26 27
2 29 23 3d0046 1 32 8 0 0 #STATE_DATA
2 30 23 300039 1 32 8 0 0 #STATE_TAIL
2 31 23 1f0039 2 1a 20208 29 30 32 0 aa aa 10aa 1aa aa aa aa aa
2 32 23 28002b 2 1 1c 0 0 tail
2 33 23 200024 1 1 18 0 0 valid
2 34 23 20002b 2 8 2033c 32 33 1 0 102
2 35 23 1f0046 2 19 202b8 31 34 16 0 aa aa 10aa 1aa
2 36 23 12001b 0 1 400 0 0 next_state
2 37 23 120046 2 37 602a 35 36
2 38 24 3d0046 1 32 8 0 0 #STATE_IDLE
2 39 24 300039 1 32 8 0 0 #STATE_HEAD
2 40 24 1f0039 2 1a 20208 38 39 32 0 1aa 10aa aa aa aa aa aa aa
2 41 24 28002b 2 1 c 0 0 head
2 42 24 200024 2 1 c 0 0 valid
2 43 24 20002b 2 8 2024c 41 42 1 0 1002
2 44 24 1f0046 2 19 20288 40 43 16 0 1aa 10aa aa aa
2 45 24 12001b 0 1 400 0 0 next_state
2 46 24 120046 2 37 600a 44 45
2 47 24 5000e 1 32 8 0 0 #STATE_TAIL
2 48 20 9000d 19 1 a 0 0 state
2 49 24 0 3 2d 2420e 47 48 1 0 102
2 50 23 5000e 1 32 8 0 0 #STATE_DATA
2 51 23 0 5 2d 2020e 50 48 1 0 1102
2 52 22 5000e 1 32 8 0 0 #STATE_HEAD
2 53 22 0 7 2d 2020e 52 48 1 0 1102
2 54 21 5000e 1 32 8 0 0 #STATE_IDLE
2 55 21 0 a 2d 2020e 54 48 1 0 1102
2 56 18 230026 5 1 c 0 0 tail
2 57 18 230026 0 2a 20000 0 0 2 0 110a
2 58 18 230026 5 29 20008 56 57 1 0 2
2 59 18 1a001e 3 1 c 0 0 valid
2 60 18 1a001e 0 2a 20000 0 0 2 0 110a
2 61 18 1a001e 3 29 20008 59 60 1 0 2
2 62 18 120015 5 1 c 0 0 head
2 63 18 120015 0 2a 20000 0 0 2 0 110a
2 64 18 120015 5 29 20008 62 63 1 0 2
2 65 18 9000d 8 1 8 0 0 state
2 66 18 9000d 0 2a 20000 0 0 17 0 11aa 11aa 11aa 11aa 2
2 67 18 9000d 8 29 20008 65 66 1 0 2
2 68 18 90015 9 2b 20008 64 67 1 0 2
2 69 18 9001e 9 2b 20008 61 68 1 0 2
2 70 18 90026 15 2b 2100a 58 69 1 0 2
2 71 60 7000a 1 0 20004 0 0 1 1 0
2 72 60 10003 0 1 400 0 0 clk
2 73 60 1000a 1 37 1006 71 72
2 74 61 1c001e 31 1 1c 0 0 clk
2 75 61 1b001b 31 1b 2002c 74 0 1 0 1102
2 76 61 150017 0 1 400 0 0 clk
2 77 61 15001e 31 37 602e 75 76
2 78 61 120012 1 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 79 61 120012 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 80 61 100013 63 2c 2000a 78 79 32 0 aa aa aa aa aa aa aa aa
2 81 0 0 9 1 f00a 0 0 next_state
2 82 0 0 8 1 f00a 0 0 state
1 #STATE_IDLE 0 0 0 32 0 1 0 0 0 0 0 0 0
1 #STATE_HEAD 0 0 0 32 0 0 1 0 0 0 0 0 0
1 #STATE_DATA 0 0 0 32 0 0 0 1 0 0 0 0 0
1 #STATE_TAIL 0 0 0 32 0 0 0 0 1 0 0 0 0
1 clk 0 8 3000c 1 16 1102
1 reset 0 9 3000c 1 0 1002
1 head 0 10 3000c 1 0 1102
1 tail 0 11 3000c 1 0 1102
1 valid 0 12 3000c 1 0 1102
1 state 0 13 3000c 16 0 11aa 11aa 11aa 11aa
1 next_state 0 14 3000c 16 16 11aa 11aa 11aa 11aa
4 82 82 82
4 81 81 81
4 7 10 10
4 10 7 0
4 46 70 70
4 49 46 70
4 37 70 70
4 51 37 49
4 28 70 70
4 53 28 51
4 19 70 70
4 55 19 53
4 70 55 0
4 77 80 80
4 80 77 0
4 73 80 80
6 82 81 1 10,10,08,,21,20,,010220,,0120,02,0120,20,01,0220,0102,,0201,0202,21,,,02
*/

/* OUTPUT fsm3.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm3.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm3.v                     9/    0/    9      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm3.v                    12/   25/   37       32%            13/   24/   37       35%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      state                     0->1: 16'h1111
      ......................... 1->0: 16'h1111 ...
      next_state                0->1: 16'h1111
      ......................... 1->0: 16'h1111 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm3.v                             23/  14/  37       62%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    state <= reset ? STATE_IDLE : next_state
                             |--------------1--------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    case( state ) 
                          |-1-|   
                    STATE_IDLE :

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm3.v                    4/  ? /  ?        ? %            8/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          16'h0001
          16'h0010
          16'h0100
          16'h1000

        Hit State Transitions

          From State    To State  
          ==========    ==========
          16'h0001   -> 16'h0001  
          16'h0001   -> 16'h0010  
          16'h0010   -> 16'h0100  
          16'h0100   -> 16'h0100  
          16'h0100   -> 16'h1000  
          16'h1000   -> 16'h0010  
          16'h0010   -> 16'h1000  
          16'h1000   -> 16'h0001  



*/

/* OUTPUT fsm3.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm3.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm3.v                     9/    0/    9      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm3.v                    12/   25/   37       32%            13/   24/   37       35%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      state                     0->1: 16'h1111
      ......................... 1->0: 16'h1111 ...
      next_state                0->1: 16'h1111
      ......................... 1->0: 16'h1111 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm3.v                             23/  14/  37       62%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    state <= reset ? STATE_IDLE : next_state
                             |--------------1--------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    case( state ) STATE_IDLE :
                          |-1-|               

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm3.v                    4/  ? /  ?        ? %            8/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          16'h0001
          16'h0010
          16'h0100
          16'h1000

        Hit State Transitions

          From State    To State  
          ==========    ==========
          16'h0001   -> 16'h0001  
          16'h0001   -> 16'h0010  
          16'h0010   -> 16'h0100  
          16'h0100   -> 16'h0100  
          16'h0100   -> 16'h1000  
          16'h1000   -> 16'h0010  
          16'h0010   -> 16'h1000  
          16'h1000   -> 16'h0001  



*/

/* OUTPUT fsm3.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm3.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    0/    9      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         12/   25/   37       32%            13/   24/   37       35%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      state                     0->1: 16'h1111
      ......................... 1->0: 16'h1111 ...
      next_state                0->1: 16'h1111
      ......................... 1->0: 16'h1111 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            23/  14/  37       62%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    state <= reset ? STATE_IDLE : next_state
                             |--------------1--------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    case( state ) 
                          |-1-|   
                    STATE_IDLE :

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         4/  ? /  ?        ? %            8/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          16'h0001
          16'h0010
          16'h0100
          16'h1000

        Hit State Transitions

          From State    To State  
          ==========    ==========
          16'h0001   -> 16'h0001  
          16'h0001   -> 16'h0010  
          16'h0010   -> 16'h0100  
          16'h0100   -> 16'h0100  
          16'h0100   -> 16'h1000  
          16'h1000   -> 16'h0010  
          16'h0010   -> 16'h1000  
          16'h1000   -> 16'h0001  



*/

/* OUTPUT fsm3.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm3.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    0/    9      100%


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         12/   25/   37       32%            13/   24/   37       35%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...
      state                     0->1: 16'h1111
      ......................... 1->0: 16'h1111 ...
      next_state                0->1: 16'h1111
      ......................... 1->0: 16'h1111 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            23/  14/  37       62%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             16:    state <= reset ? STATE_IDLE : next_state
                             |--------------1--------------|

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    case( state ) STATE_IDLE :
                          |-1-|               

        Expression 1   (1/2)
        ^^^^^^^^^^^^^ - 
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             21:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & tail) ? STATE_TAIL : STATE_DATA
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *          

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & head) ? STATE_HEAD : STATE_IDLE
                                 |-----1------|                          
                                 |------------------2-------------------|

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         4/  ? /  ?        ? %            8/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm3.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state)

        Hit States

          States
          ======
          16'h0001
          16'h0010
          16'h0100
          16'h1000

        Hit State Transitions

          From State    To State  
          ==========    ==========
          16'h0001   -> 16'h0001  
          16'h0001   -> 16'h0010  
          16'h0010   -> 16'h0100  
          16'h0100   -> 16'h0100  
          16'h0100   -> 16'h1000  
          16'h1000   -> 16'h0010  
          16'h0010   -> 16'h1000  
          16'h1000   -> 16'h0001  



*/
