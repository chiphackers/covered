module main;

parameter [1:0] STATE_IDLE = 2'b00,
                STATE_HEAD = 2'b01,
                STATE_DATA = 2'b10,
	        STATE_TAIL = 2'b11;

reg            clock;
reg            reset;
reg  [1:0]     state;
reg  [2:0]     next_state;
wire           msg_ip;
reg            head;
reg            tail;
reg            valid;

always @(posedge clock) state <= reset ? {1'b0,STATE_IDLE} : next_state;

always @(state or head or valid or tail)
  begin
   case( state )
     STATE_IDLE:  next_state = (valid & head) ? {1'b1,STATE_HEAD} : {1'b0,STATE_IDLE};
     STATE_HEAD:  next_state = (valid & tail) ? {1'b1,STATE_TAIL} : {1'b1,STATE_DATA};
     STATE_DATA:  next_state = (valid & tail) ? {1'b1,STATE_TAIL} : {1'b1,STATE_DATA};
     STATE_TAIL:  next_state = (valid & head) ? {1'b1,STATE_HEAD} : {1'b0,STATE_IDLE};
   endcase
  end

assign msg_ip = next_state[2];

initial begin
	$dumpfile( "fsm5.vcd" );
	$dumpvars( 0, main );
	reset = 1'b1;
	valid = 1'b0;
	head  = 1'b0;
	tail  = 1'b0;
	#20;
	reset = 1'b0;
	@(posedge clock);
        head  <= 1'b1;
        valid <= 1'b1;
	@(posedge clock);
	head  <= 1'b0;
	tail  <= 1'b1;
	@(posedge clock);
	tail  <= 1'b0;
	valid <= 1'b0;
	#20;
	$finish;
end

initial begin
	clock = 1'b0;
	forever #(1) clock = ~clock;
end

endmodule

/* HEADER
GROUPS fsm5 all iv vcs vcd lxt
SIM    fsm5 all iv vcd  : iverilog fsm5.v; ./a.out                             : fsm5.vcd
SIM    fsm5 all iv lxt  : iverilog fsm5.v; ./a.out -lxt2; mv fsm5.vcd fsm5.lxt : fsm5.lxt
SIM    fsm5 all vcs vcd : vcs fsm5.v; ./simv                                   : fsm5.vcd
SCORE  fsm5.vcd     : -t main -vcd fsm5.vcd -o fsm5.cdd -y lib -v fsm5.v -F main=state,next_state[1:0] : fsm5.cdd
SCORE  fsm5.lxt     : -t main -lxt fsm5.lxt -o fsm5.cdd -y lib -v fsm5.v -F main=state,next_state[1:0] : fsm5.cdd
REPORT fsm5.cdd 1   : -d v -o fsm5.rptM fsm5.cdd                         : fsm5.rptM
REPORT fsm5.cdd 2   : -d v -w -o fsm5.rptWM fsm5.cdd                     : fsm5.rptWM
REPORT fsm5.cdd 3   : -d v -i -o fsm5.rptI fsm5.cdd                      : fsm5.rptI
REPORT fsm5.cdd 4   : -d v -w -i -o fsm5.rptWI fsm5.cdd                  : fsm5.rptWI
*/

/* OUTPUT fsm5.cdd
5 1 * 6 0 0 0 0
3 0 main main fsm5.v 1 58
2 1 17 3d0046 5 1 c 0 0 next_state
2 2 17 2f0038 1 32 4 0 0 #STATE_IDLE
2 3 17 2a002d 1 0 20004 0 0 1 1 0
2 4 17 2a0038 1 31 20044 2 3 3 0 2a
2 5 17 290039 1 26 20004 4 0 3 0 2a
2 6 17 210039 7 1a 200cc 1 5 3 0 772a
2 7 17 210025 2 1 c 0 0 reset
2 8 17 210046 7 19 201cc 6 7 2 0 330a
2 9 17 18001c 0 1 400 0 0 state
2 10 17 180046 17 38 600e 8 9
2 11 17 110015 2e 1 c 0 0 clock
2 12 17 9000f 0 2a 20000 0 0 2 0 a
2 13 17 90015 46 27 2100a 11 12 1 0 2
2 14 22 4a0053 1 32 4 0 0 #STATE_IDLE
2 15 22 450048 1 0 20004 0 0 1 1 0
2 16 22 450053 1 31 20044 14 15 3 0 2a
2 17 22 440054 1 26 20004 16 0 3 0 2a
2 18 22 36003f 1 32 8 0 0 #STATE_HEAD
2 19 22 310034 1 0 20008 0 0 1 1 1
2 20 22 31003f 1 31 20208 18 19 3 0 2a
2 21 22 300040 1 26 20008 20 0 3 0 2a
2 22 22 1f0040 3 1a 2010c 17 21 3 0 552a
2 23 22 28002b 3 1 c 0 0 head
2 24 22 200024 3 1 c 0 0 valid
2 25 22 20002b 3 8 2024c 23 24 1 0 1102
2 26 22 1f0054 3 19 2024c 22 25 3 0 552a
2 27 22 12001b 0 1 400 0 0 next_state
2 28 22 120054 3 37 600e 26 27
2 29 23 4a0053 1 32 8 0 0 #STATE_DATA
2 30 23 450048 1 0 20008 0 0 1 1 1
2 31 23 450053 1 31 20208 29 30 3 0 2a
2 32 23 440054 1 26 20008 31 0 3 0 2a
2 33 23 36003f 1 32 8 0 0 #STATE_TAIL
2 34 23 310034 1 0 20008 0 0 1 1 1
2 35 23 31003f 1 31 20208 33 34 3 0 2a
2 36 23 300040 1 26 20008 35 0 3 0 2a
2 37 23 1f0040 1 1a 20208 32 36 3 0 2a
2 38 23 28002b 1 1 18 0 0 tail
2 39 23 200024 1 1 18 0 0 valid
2 40 23 20002b 1 8 20238 38 39 1 0 2
2 41 23 1f0054 1 19 20238 37 40 3 0 2a
2 42 23 12001b 0 1 400 0 0 next_state
2 43 23 120054 1 37 602a 41 42
2 44 24 4a0053 0 32 10 0 0 #STATE_DATA
2 45 24 450048 0 0 20010 0 0 1 1 1
2 46 24 450053 0 31 20030 44 45 3 0 2a
2 47 24 440054 0 26 20020 46 0 3 0 2a
2 48 24 36003f 0 32 10 0 0 #STATE_TAIL
2 49 24 310034 0 0 20010 0 0 1 1 1
2 50 24 31003f 0 31 20030 48 49 3 0 2a
2 51 24 300040 0 26 20020 50 0 3 0 2a
2 52 24 1f0040 0 1a 20030 47 51 3 0 2a
2 53 24 28002b 0 1 10 0 0 tail
2 54 24 200024 0 1 10 0 0 valid
2 55 24 20002b 0 8 20030 53 54 1 0 2
2 56 24 1f0054 0 19 20030 52 55 3 0 2a
2 57 24 12001b 0 1 400 0 0 next_state
2 58 24 120054 0 37 6022 56 57
2 59 25 4a0053 1 32 4 0 0 #STATE_IDLE
2 60 25 450048 1 0 20004 0 0 1 1 0
2 61 25 450053 1 31 20044 59 60 3 0 2a
2 62 25 440054 1 26 20004 61 0 3 0 2a
2 63 25 36003f 1 32 8 0 0 #STATE_HEAD
2 64 25 310034 1 0 20008 0 0 1 1 1
2 65 25 31003f 1 31 20208 63 64 3 0 2a
2 66 25 300040 1 26 20008 65 0 3 0 2a
2 67 25 1f0040 1 1a 20104 62 66 3 0 2a
2 68 25 28002b 1 1 4 0 0 head
2 69 25 200024 1 1 4 0 0 valid
2 70 25 20002b 1 8 20044 68 69 1 0 2
2 71 25 1f0054 1 19 20044 67 70 3 0 2a
2 72 25 12001b 0 1 400 0 0 next_state
2 73 25 120054 1 37 6006 71 72
2 74 25 5000e 1 32 8 0 0 #STATE_TAIL
2 75 21 9000d d 1 e 0 0 state
2 76 25 0 2 2d 2420e 74 75 1 0 102
2 77 24 5000e 1 32 8 0 0 #STATE_DATA
2 78 24 0 2 2d 20206 77 75 1 0 2
2 79 23 5000e 1 32 8 0 0 #STATE_HEAD
2 80 23 0 3 2d 2020e 79 75 1 0 1102
2 81 22 5000e 1 32 4 0 0 #STATE_IDLE
2 82 22 0 6 2d 2014e 81 75 1 0 1102
2 83 19 230026 3 1 c 0 0 tail
2 84 19 230026 0 2a 20000 0 0 2 0 110a
2 85 19 230026 3 29 20008 83 84 1 0 2
2 86 19 1a001e 3 1 c 0 0 valid
2 87 19 1a001e 0 2a 20000 0 0 2 0 110a
2 88 19 1a001e 3 29 20008 86 87 1 0 2
2 89 19 120015 3 1 c 0 0 head
2 90 19 120015 0 2a 20000 0 0 2 0 110a
2 91 19 120015 3 29 20008 89 90 1 0 2
2 92 19 9000d 5 1 c 0 0 state
2 93 19 9000d 0 2a 20000 0 0 3 0 332a
2 94 19 9000d 5 29 20008 92 93 1 0 2
2 95 19 90015 6 2b 20008 91 94 1 0 2
2 96 19 9001e 6 2b 20008 88 95 1 0 2
2 97 19 90026 d 2b 2100a 85 96 1 0 2
2 98 29 1b001b 6 0 20008 0 0 32 64 4 0 0 0 0 0 0 0
2 99 29 10001c 6 23 c 0 98 next_state
2 100 29 7000c 0 1 400 0 0 msg_ip
2 101 29 7001c 6 35 f00e 99 100
2 102 54 9000c 1 0 20004 0 0 1 1 0
2 103 54 10005 0 1 400 0 0 clock
2 104 54 1000c 1 37 1006 102 103
2 105 55 17001b 2d 1 1c 0 0 clock
2 106 55 160016 2d 1b 2002c 105 0 1 0 1102
2 107 55 e0012 0 1 400 0 0 clock
2 108 55 e001b 2d 37 602e 106 107
2 109 55 b000b 1 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 110 55 b000b 1 0 20008 0 0 32 64 55 55 55 55 55 55 55 55
2 111 55 9000c 5b 2c 2000a 109 110 32 0 aa aa aa aa aa aa aa aa
2 112 0 0 1 0 20004 0 0 32 64 0 0 0 0 0 0 0 0
2 113 0 0 6 0 20008 0 0 32 64 1 0 0 0 0 0 0 0
2 114 0 0 6 24 f10e 112 113 next_state
2 115 0 0 5 1 f00e 0 0 state
1 #STATE_IDLE 0 0 0 2 0 0
1 #STATE_HEAD 0 0 0 2 0 1
1 #STATE_DATA 0 0 0 2 0 4
1 #STATE_TAIL 0 0 0 2 0 5
1 clock 0 8 3000f 1 16 1102
1 reset 0 9 3000f 1 0 1002
1 state 0 10 3000f 2 0 330a
1 next_state 0 11 3000f 3 16 772a
1 msg_ip 0 12 3000f 1 0 1102
1 head 0 13 3000f 1 0 1102
1 tail 0 14 3000f 1 0 1102
1 valid 0 15 3000f 1 0 1102
4 115 115 115
4 114 114 114
4 10 13 13
4 13 10 0
4 73 97 97
4 76 73 97
4 58 97 97
4 78 58 76
4 43 97 97
4 80 43 78
4 28 97 97
4 82 28 80
4 97 82 0
4 101 101 101
4 108 111 111
4 111 108 0
4 104 111 111
6 115 114 1 02,04,04,,01,21,e1,8101
*/

/* OUTPUT fsm5.rptM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm5.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.v                     9/    1/   10       90%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           24:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.v                    10/    1/   11       91%            11/    0/   11      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm5.v                             41/  16/  57       72%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:    next_state = (valid & head) ? {1'b1, STATE_HEAD} : {1'b0, STATE_IDLE}
                                 |-----1------|                                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & head) ? {1'b1, STATE_HEAD} : {1'b0, STATE_IDLE}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.v                    3/  ? /  ?        ? %            4/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state[1:0])

        Hit States

          States
          ======
          2'h0
          2'h1
          2'h3

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      
          2'h0       -> 2'h1      
          2'h1       -> 2'h3      
          2'h3       -> 2'h0      



*/

/* OUTPUT fsm5.rptWM
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm5.cdd

* Reported by                    : Module

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                 Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.v                     9/    1/   10       90%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           24:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function      Filename                         Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.v                    10/    1/   11       91%            11/    0/   11      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Module/Task/Function                Filename                                Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                              fsm5.v                             41/  16/  57       72%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:    next_state = (valid & head) ? {1'b1, STATE_HEAD} : {1'b0, STATE_IDLE}
                                 |-----1------|                                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & head) ? {1'b1, STATE_HEAD} : {1'b0, STATE_IDLE}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Module/Task/Function      Filename                Hit/Miss/Total    Percent Hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  main                    fsm5.v                    3/  ? /  ?        ? %            4/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state[1:0])

        Hit States

          States
          ======
          2'h0
          2'h1
          2'h3

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      
          2'h0       -> 2'h1      
          2'h1       -> 2'h3      
          2'h3       -> 2'h0      



*/

/* OUTPUT fsm5.rptI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm5.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    1/   10       90%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           24:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         10/    1/   11       91%            11/    0/   11      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            41/  16/  57       72%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:    next_state = (valid & head) ? {1'b1, STATE_HEAD} : {1'b0, STATE_IDLE}
                                 |-----1------|                                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & head) ? {1'b1, STATE_HEAD} : {1'b0, STATE_IDLE}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         3/  ? /  ?        ? %            4/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state[1:0])

        Hit States

          States
          ======
          2'h0
          2'h1
          2'h3

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      
          2'h0       -> 2'h1      
          2'h1       -> 2'h3      
          2'h3       -> 2'h0      



*/

/* OUTPUT fsm5.rptWI
                             ::::::::::::::::::::::::::::::::::::::::::::::::::
                             ::                                              ::
                             ::  Covered -- Verilog Coverage Verbose Report  ::
                             ::                                              ::
                             ::::::::::::::::::::::::::::::::::::::::::::::::::


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   GENERAL INFORMATION   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
* Report generated from CDD file : fsm5.cdd

* Reported by                    : Instance

~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   LINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                           Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                          9/    1/   10       90%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Lines

           24:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   TOGGLE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                   Toggle 0 -> 1                       Toggle 1 -> 0
                                                   Hit/ Miss/Total    Percent hit      Hit/ Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         10/    1/   11       91%            11/    0/   11      100%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Signals not getting 100% toggle coverage

      Signal                    Toggle
      ---------------------------------------------------------------------------------------------------------
      reset                     0->1: 1'h0
      ......................... 1->0: 1'h1 ...


~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   COMBINATIONAL LOGIC COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
Instance                                                                    Logic Combinations
                                                                      Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                                            41/  16/  57       72%
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
    Missed Combinations  (* = missed value)

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             22:    next_state = (valid & head) ? {1'b1, STATE_HEAD} : {1'b0, STATE_IDLE}
                                 |-----1------|                                          

        Expression 1   (2/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *     

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             23:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *     

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *    

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             24:    next_state = (valid & tail) ? {1'b1, STATE_TAIL} : {1'b1, STATE_DATA}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (0/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
         *    *    *    *

        Expression 2   (0/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
         *   *

      =========================================================================================================
       Line #     Expression
      =========================================================================================================
             25:    next_state = (valid & head) ? {1'b1, STATE_HEAD} : {1'b0, STATE_IDLE}
                                 |-----1------|                                          
                                 |--------------------------2---------------------------|

        Expression 1   (1/4)
        ^^^^^^^^^^^^^ - &
         LR | LR | LR | LR 
        =00=|=01=|=10=|=11=
              *    *    *

        Expression 2   (1/2)
        ^^^^^^^^^^^^^ - ?:
         E | E
        =0=|=1=
             *



~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~   FINITE STATE MACHINE COVERAGE RESULTS   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
                                                               State                             Arc
Instance                                          Hit/Miss/Total    Percent hit    Hit/Miss/Total    Percent hit
---------------------------------------------------------------------------------------------------------------------
  <NA>.main                                         3/  ? /  ?        ? %            4/  ? /  ?        ? %
---------------------------------------------------------------------------------------------------------------------

    Module: main, File: fsm5.v, Instance: <NA>.main
    -------------------------------------------------------------------------------------------------------------
      FSM input state (state), output state (next_state[1:0])

        Hit States

          States
          ======
          2'h0
          2'h1
          2'h3

        Hit State Transitions

          From State    To State  
          ==========    ==========
          2'h0       -> 2'h0      
          2'h0       -> 2'h1      
          2'h1       -> 2'h3      
          2'h3       -> 2'h0      



*/
